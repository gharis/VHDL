
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sin_inv is
port
(
   clk               :  IN  std_logic;
	reset 				: 	IN STD_LOGIC;
	clk_50				: 	IN STD_LOGIC;
	avs_s0_address		: 	IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	avs_s0_read			: 	IN STD_LOGIC;
	avs_s0_write		: 	IN STD_LOGIC;
	avs_s0_readdata	: 	OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
	avs_s0_writedata	: 	IN STD_LOGIC_VECTOR(31 DOWNTO 0)
);
end sin_inv;


architecture rtl of sin_inv is
    signal reset_n    : std_logic;
	 signal theta_inv     : std_logic_vector(31 downto 0);
    signal clk_en     : std_logic;
    signal sin_inv      : signed(31 downto 0);
	-- signal sin_inv_data   : signed(31 downto 0);
	 signal sin_inv_data   : integer;

	 type my_array is array (0 to 6) of std_logic_vector(2 downto 0);
	 signal sequence: my_array;
   
	 type t_Integer_Array is array (0 to 3) of integer; --4 elements
	
	 type int_array is array (0 to 512) of integer; --first define the type of array.
signal led : std_logic_vector(7 downto 0); 
begin




   AV_READ: PROCESS(clk)
	BEGIN
		IF rising_edge(clk) THEN
			IF (reset='1') THEN
				avs_s0_readdata <= x"00000000";
				ELSIF (avs_s0_read='1') THEN
					IF (avs_s0_address = x"00" )THEN
						avs_s0_readdata 	<=		std_logic_vector(sin_inv(31 downto 0)) AND x"FFFFFFFF";
					ELSE avs_s0_readdata <= x"0000ffff";
				END IF;		
			END IF;
		END IF;
	END PROCESS;
		 
	  AV_WRITE: PROCESS(clk)
	  BEGIN
        IF rising_edge(clk) THEN
            IF (reset='1') THEN
                led <= "00001111";
            ELSIF (avs_s0_write='1') THEN               
					 IF (avs_s0_address = x"00" )THEN
                    theta_inv 				<= avs_s0_writedata(31 downto 0); 

					 ELSIF (avs_s0_address = x"01") THEN
                    clk_en 		   <= avs_s0_writedata(0);
						  reset_n         <= NOT(clk_en);
					 ELSE led 						<= "11110000";
					 END IF; 
            END IF;
        END IF;
	  END PROCESS;	





 SIN_inv_lookup: process(clk_50)
 variable theta_int_inv  : integer range -1000 to 1000 := 0;

 begin
   if(reset_n = '1')then
       sin_inv <= to_signed(3000,32); 
   elsif(rising_edge(clk_50)) then
      if clk_en = '1' then
		theta_int_inv := to_integer(signed(theta_inv));
      --sin_inv <=  sin_inv_data;

      sin_inv <=  to_signed(sin_inv_data,32);
--
--      case theta_int_inv is
--			when -1000 => sin_inv_data <= to_signed(-90,32);
--			when -999 => sin_inv_data <= to_signed(-87,32);
--			when -998 => sin_inv_data <= to_signed(-86,32);
--			when -997 => sin_inv_data <= to_signed(-86,32);
--			when -996 => sin_inv_data <= to_signed(-85,32);
--			when -995 => sin_inv_data <= to_signed(-84,32);
--			when -994 => sin_inv_data <= to_signed(-84,32);
--			when -993 => sin_inv_data <= to_signed(-83,32);
--			when -992 => sin_inv_data <= to_signed(-83,32);
--			when -991 => sin_inv_data <= to_signed(-82,32);
--			when -990 => sin_inv_data <= to_signed(-82,32);
--			when -989 => sin_inv_data <= to_signed(-81,32);
--			when -988 => sin_inv_data <= to_signed(-81,32);
--			when -987 => sin_inv_data <= to_signed(-81,32);
--			when -986 => sin_inv_data <= to_signed(-80,32);
--			when -985 => sin_inv_data <= to_signed(-80,32);
--			when -984 => sin_inv_data <= to_signed(-80,32);
--			when -983 => sin_inv_data <= to_signed(-79,32);
--			when -982 => sin_inv_data <= to_signed(-79,32);
--			when -981 => sin_inv_data <= to_signed(-79,32);
--			when -980 => sin_inv_data <= to_signed(-79,32);
--			when -979 => sin_inv_data <= to_signed(-78,32);
--			when -978 => sin_inv_data <= to_signed(-78,32);
--			when -977 => sin_inv_data <= to_signed(-78,32);
--			when -976 => sin_inv_data <= to_signed(-77,32);
--			when -975 => sin_inv_data <= to_signed(-77,32);
--			when -974 => sin_inv_data <= to_signed(-77,32);
--			when -973 => sin_inv_data <= to_signed(-77,32);
--			when -972 => sin_inv_data <= to_signed(-76,32);
--			when -971 => sin_inv_data <= to_signed(-76,32);
--			when -970 => sin_inv_data <= to_signed(-76,32);
--			when -969 => sin_inv_data <= to_signed(-76,32);
--			when -968 => sin_inv_data <= to_signed(-75,32);
--			when -967 => sin_inv_data <= to_signed(-75,32);
--			when -966 => sin_inv_data <= to_signed(-75,32);
--			when -965 => sin_inv_data <= to_signed(-75,32);
--			when -964 => sin_inv_data <= to_signed(-75,32);
--			when -963 => sin_inv_data <= to_signed(-74,32);
--			when -962 => sin_inv_data <= to_signed(-74,32);
--			when -961 => sin_inv_data <= to_signed(-74,32);
--			when -960 => sin_inv_data <= to_signed(-74,32);
--			when -959 => sin_inv_data <= to_signed(-74,32);
--			when -958 => sin_inv_data <= to_signed(-73,32);
--			when -957 => sin_inv_data <= to_signed(-73,32);
--			when -956 => sin_inv_data <= to_signed(-73,32);
--			when -955 => sin_inv_data <= to_signed(-73,32);
--			when -954 => sin_inv_data <= to_signed(-73,32);
--			when -953 => sin_inv_data <= to_signed(-72,32);
--			when -952 => sin_inv_data <= to_signed(-72,32);
--			when -951 => sin_inv_data <= to_signed(-72,32);
--			when -950 => sin_inv_data <= to_signed(-72,32);
--			when -949 => sin_inv_data <= to_signed(-72,32);
--			when -948 => sin_inv_data <= to_signed(-71,32);
--			when -947 => sin_inv_data <= to_signed(-71,32);
--			when -946 => sin_inv_data <= to_signed(-71,32);
--			when -945 => sin_inv_data <= to_signed(-71,32);
--			when -944 => sin_inv_data <= to_signed(-71,32);
--			when -943 => sin_inv_data <= to_signed(-71,32);
--			when -942 => sin_inv_data <= to_signed(-70,32);
--			when -941 => sin_inv_data <= to_signed(-70,32);
--			when -940 => sin_inv_data <= to_signed(-70,32);
--			when -939 => sin_inv_data <= to_signed(-70,32);
--			when -938 => sin_inv_data <= to_signed(-70,32);
--			when -937 => sin_inv_data <= to_signed(-70,32);
--			when -936 => sin_inv_data <= to_signed(-69,32);
--			when -935 => sin_inv_data <= to_signed(-69,32);
--			when -934 => sin_inv_data <= to_signed(-69,32);
--			when -933 => sin_inv_data <= to_signed(-69,32);
--			when -932 => sin_inv_data <= to_signed(-69,32);
--			when -931 => sin_inv_data <= to_signed(-69,32);
--			when -930 => sin_inv_data <= to_signed(-68,32);
--			when -929 => sin_inv_data <= to_signed(-68,32);
--			when -928 => sin_inv_data <= to_signed(-68,32);
--			when -927 => sin_inv_data <= to_signed(-68,32);
--			when -926 => sin_inv_data <= to_signed(-68,32);
--			when -925 => sin_inv_data <= to_signed(-68,32);
--			when -924 => sin_inv_data <= to_signed(-68,32);
--			when -923 => sin_inv_data <= to_signed(-67,32);
--			when -922 => sin_inv_data <= to_signed(-67,32);
--			when -921 => sin_inv_data <= to_signed(-67,32);
--			when -920 => sin_inv_data <= to_signed(-67,32);
--			when -919 => sin_inv_data <= to_signed(-67,32);
--			when -918 => sin_inv_data <= to_signed(-67,32);
--			when -917 => sin_inv_data <= to_signed(-66,32);
--			when -916 => sin_inv_data <= to_signed(-66,32);
--			when -915 => sin_inv_data <= to_signed(-66,32);
--			when -914 => sin_inv_data <= to_signed(-66,32);
--			when -913 => sin_inv_data <= to_signed(-66,32);
--			when -912 => sin_inv_data <= to_signed(-66,32);
--			when -911 => sin_inv_data <= to_signed(-66,32);
--			when -910 => sin_inv_data <= to_signed(-66,32);
--			when -909 => sin_inv_data <= to_signed(-65,32);
--			when -908 => sin_inv_data <= to_signed(-65,32);
--			when -907 => sin_inv_data <= to_signed(-65,32);
--			when -906 => sin_inv_data <= to_signed(-65,32);
--			when -905 => sin_inv_data <= to_signed(-65,32);
--			when -904 => sin_inv_data <= to_signed(-65,32);
--			when -903 => sin_inv_data <= to_signed(-65,32);
--			when -902 => sin_inv_data <= to_signed(-64,32);
--			when -901 => sin_inv_data <= to_signed(-64,32);
--			when -900 => sin_inv_data <= to_signed(-64,32);
--			when -899 => sin_inv_data <= to_signed(-64,32);
--			when -898 => sin_inv_data <= to_signed(-64,32);
--			when -897 => sin_inv_data <= to_signed(-64,32);
--			when -896 => sin_inv_data <= to_signed(-64,32);
--			when -895 => sin_inv_data <= to_signed(-64,32);
--			when -894 => sin_inv_data <= to_signed(-63,32);
--			when -893 => sin_inv_data <= to_signed(-63,32);
--			when -892 => sin_inv_data <= to_signed(-63,32);
--			when -891 => sin_inv_data <= to_signed(-63,32);
--			when -890 => sin_inv_data <= to_signed(-63,32);
--			when -889 => sin_inv_data <= to_signed(-63,32);
--			when -888 => sin_inv_data <= to_signed(-63,32);
--			when -887 => sin_inv_data <= to_signed(-62,32);
--			when -886 => sin_inv_data <= to_signed(-62,32);
--			when -885 => sin_inv_data <= to_signed(-62,32);
--			when -884 => sin_inv_data <= to_signed(-62,32);
--			when -883 => sin_inv_data <= to_signed(-62,32);
--			when -882 => sin_inv_data <= to_signed(-62,32);
--			when -881 => sin_inv_data <= to_signed(-62,32);
--			when -880 => sin_inv_data <= to_signed(-62,32);
--			when -879 => sin_inv_data <= to_signed(-62,32);
--			when -878 => sin_inv_data <= to_signed(-61,32);
--			when -877 => sin_inv_data <= to_signed(-61,32);
--			when -876 => sin_inv_data <= to_signed(-61,32);
--			when -875 => sin_inv_data <= to_signed(-61,32);
--			when -874 => sin_inv_data <= to_signed(-61,32);
--			when -873 => sin_inv_data <= to_signed(-61,32);
--			when -872 => sin_inv_data <= to_signed(-61,32);
--			when -871 => sin_inv_data <= to_signed(-61,32);
--			when -870 => sin_inv_data <= to_signed(-60,32);
--			when -869 => sin_inv_data <= to_signed(-60,32);
--			when -868 => sin_inv_data <= to_signed(-60,32);
--			when -867 => sin_inv_data <= to_signed(-60,32);
--			when -866 => sin_inv_data <= to_signed(-60,32);
--			when -865 => sin_inv_data <= to_signed(-60,32);
--			when -864 => sin_inv_data <= to_signed(-60,32);
--			when -863 => sin_inv_data <= to_signed(-60,32);
--			when -862 => sin_inv_data <= to_signed(-60,32);
--			when -861 => sin_inv_data <= to_signed(-59,32);
--			when -860 => sin_inv_data <= to_signed(-59,32);
--			when -859 => sin_inv_data <= to_signed(-59,32);
--			when -858 => sin_inv_data <= to_signed(-59,32);
--			when -857 => sin_inv_data <= to_signed(-59,32);
--			when -856 => sin_inv_data <= to_signed(-59,32);
--			when -855 => sin_inv_data <= to_signed(-59,32);
--			when -854 => sin_inv_data <= to_signed(-59,32);
--			when -853 => sin_inv_data <= to_signed(-59,32);
--			when -852 => sin_inv_data <= to_signed(-58,32);
--			when -851 => sin_inv_data <= to_signed(-58,32);
--			when -850 => sin_inv_data <= to_signed(-58,32);
--			when -849 => sin_inv_data <= to_signed(-58,32);
--			when -848 => sin_inv_data <= to_signed(-58,32);
--			when -847 => sin_inv_data <= to_signed(-58,32);
--			when -846 => sin_inv_data <= to_signed(-58,32);
--			when -845 => sin_inv_data <= to_signed(-58,32);
--			when -844 => sin_inv_data <= to_signed(-58,32);
--			when -843 => sin_inv_data <= to_signed(-57,32);
--			when -842 => sin_inv_data <= to_signed(-57,32);
--			when -841 => sin_inv_data <= to_signed(-57,32);
--			when -840 => sin_inv_data <= to_signed(-57,32);
--			when -839 => sin_inv_data <= to_signed(-57,32);
--			when -838 => sin_inv_data <= to_signed(-57,32);
--			when -837 => sin_inv_data <= to_signed(-57,32);
--			when -836 => sin_inv_data <= to_signed(-57,32);
--			when -835 => sin_inv_data <= to_signed(-57,32);
--			when -834 => sin_inv_data <= to_signed(-57,32);
--			when -833 => sin_inv_data <= to_signed(-56,32);
--			when -832 => sin_inv_data <= to_signed(-56,32);
--			when -831 => sin_inv_data <= to_signed(-56,32);
--			when -830 => sin_inv_data <= to_signed(-56,32);
--			when -829 => sin_inv_data <= to_signed(-56,32);
--			when -828 => sin_inv_data <= to_signed(-56,32);
--			when -827 => sin_inv_data <= to_signed(-56,32);
--			when -826 => sin_inv_data <= to_signed(-56,32);
--			when -825 => sin_inv_data <= to_signed(-56,32);
--			when -824 => sin_inv_data <= to_signed(-55,32);
--			when -823 => sin_inv_data <= to_signed(-55,32);
--			when -822 => sin_inv_data <= to_signed(-55,32);
--			when -821 => sin_inv_data <= to_signed(-55,32);
--			when -820 => sin_inv_data <= to_signed(-55,32);
--			when -819 => sin_inv_data <= to_signed(-55,32);
--			when -818 => sin_inv_data <= to_signed(-55,32);
--			when -817 => sin_inv_data <= to_signed(-55,32);
--			when -816 => sin_inv_data <= to_signed(-55,32);
--			when -815 => sin_inv_data <= to_signed(-55,32);
--			when -814 => sin_inv_data <= to_signed(-54,32);
--			when -813 => sin_inv_data <= to_signed(-54,32);
--			when -812 => sin_inv_data <= to_signed(-54,32);
--			when -811 => sin_inv_data <= to_signed(-54,32);
--			when -810 => sin_inv_data <= to_signed(-54,32);
--			when -809 => sin_inv_data <= to_signed(-54,32);
--			when -808 => sin_inv_data <= to_signed(-54,32);
--			when -807 => sin_inv_data <= to_signed(-54,32);
--			when -806 => sin_inv_data <= to_signed(-54,32);
--			when -805 => sin_inv_data <= to_signed(-54,32);
--			when -804 => sin_inv_data <= to_signed(-54,32);
--			when -803 => sin_inv_data <= to_signed(-53,32);
--			when -802 => sin_inv_data <= to_signed(-53,32);
--			when -801 => sin_inv_data <= to_signed(-53,32);
--			when -800 => sin_inv_data <= to_signed(-53,32);
--			when -799 => sin_inv_data <= to_signed(-53,32);
--			when -798 => sin_inv_data <= to_signed(-53,32);
--			when -797 => sin_inv_data <= to_signed(-53,32);
--			when -796 => sin_inv_data <= to_signed(-53,32);
--			when -795 => sin_inv_data <= to_signed(-53,32);
--			when -794 => sin_inv_data <= to_signed(-53,32);
--			when -793 => sin_inv_data <= to_signed(-52,32);
--			when -792 => sin_inv_data <= to_signed(-52,32);
--			when -791 => sin_inv_data <= to_signed(-52,32);
--			when -790 => sin_inv_data <= to_signed(-52,32);
--			when -789 => sin_inv_data <= to_signed(-52,32);
--			when -788 => sin_inv_data <= to_signed(-52,32);
--			when -787 => sin_inv_data <= to_signed(-52,32);
--			when -786 => sin_inv_data <= to_signed(-52,32);
--			when -785 => sin_inv_data <= to_signed(-52,32);
--			when -784 => sin_inv_data <= to_signed(-52,32);
--			when -783 => sin_inv_data <= to_signed(-52,32);
--			when -782 => sin_inv_data <= to_signed(-51,32);
--			when -781 => sin_inv_data <= to_signed(-51,32);
--			when -780 => sin_inv_data <= to_signed(-51,32);
--			when -779 => sin_inv_data <= to_signed(-51,32);
--			when -778 => sin_inv_data <= to_signed(-51,32);
--			when -777 => sin_inv_data <= to_signed(-51,32);
--			when -776 => sin_inv_data <= to_signed(-51,32);
--			when -775 => sin_inv_data <= to_signed(-51,32);
--			when -774 => sin_inv_data <= to_signed(-51,32);
--			when -773 => sin_inv_data <= to_signed(-51,32);
--			when -772 => sin_inv_data <= to_signed(-51,32);
--			when -771 => sin_inv_data <= to_signed(-50,32);
--			when -770 => sin_inv_data <= to_signed(-50,32);
--			when -769 => sin_inv_data <= to_signed(-50,32);
--			when -768 => sin_inv_data <= to_signed(-50,32);
--			when -767 => sin_inv_data <= to_signed(-50,32);
--			when -766 => sin_inv_data <= to_signed(-50,32);
--			when -765 => sin_inv_data <= to_signed(-50,32);
--			when -764 => sin_inv_data <= to_signed(-50,32);
--			when -763 => sin_inv_data <= to_signed(-50,32);
--			when -762 => sin_inv_data <= to_signed(-50,32);
--			when -761 => sin_inv_data <= to_signed(-50,32);
--			when -760 => sin_inv_data <= to_signed(-49,32);
--			when -759 => sin_inv_data <= to_signed(-49,32);
--			when -758 => sin_inv_data <= to_signed(-49,32);
--			when -757 => sin_inv_data <= to_signed(-49,32);
--			when -756 => sin_inv_data <= to_signed(-49,32);
--			when -755 => sin_inv_data <= to_signed(-49,32);
--			when -754 => sin_inv_data <= to_signed(-49,32);
--			when -753 => sin_inv_data <= to_signed(-49,32);
--			when -752 => sin_inv_data <= to_signed(-49,32);
--			when -751 => sin_inv_data <= to_signed(-49,32);
--			when -750 => sin_inv_data <= to_signed(-49,32);
--			when -749 => sin_inv_data <= to_signed(-49,32);
--			when -748 => sin_inv_data <= to_signed(-48,32);
--			when -747 => sin_inv_data <= to_signed(-48,32);
--			when -746 => sin_inv_data <= to_signed(-48,32);
--			when -745 => sin_inv_data <= to_signed(-48,32);
--			when -744 => sin_inv_data <= to_signed(-48,32);
--			when -743 => sin_inv_data <= to_signed(-48,32);
--			when -742 => sin_inv_data <= to_signed(-48,32);
--			when -741 => sin_inv_data <= to_signed(-48,32);
--			when -740 => sin_inv_data <= to_signed(-48,32);
--			when -739 => sin_inv_data <= to_signed(-48,32);
--			when -738 => sin_inv_data <= to_signed(-48,32);
--			when -737 => sin_inv_data <= to_signed(-47,32);
--			when -736 => sin_inv_data <= to_signed(-47,32);
--			when -735 => sin_inv_data <= to_signed(-47,32);
--			when -734 => sin_inv_data <= to_signed(-47,32);
--			when -733 => sin_inv_data <= to_signed(-47,32);
--			when -732 => sin_inv_data <= to_signed(-47,32);
--			when -731 => sin_inv_data <= to_signed(-47,32);
--			when -730 => sin_inv_data <= to_signed(-47,32);
--			when -729 => sin_inv_data <= to_signed(-47,32);
--			when -728 => sin_inv_data <= to_signed(-47,32);
--			when -727 => sin_inv_data <= to_signed(-47,32);
--			when -726 => sin_inv_data <= to_signed(-47,32);
--			when -725 => sin_inv_data <= to_signed(-46,32);
--			when -724 => sin_inv_data <= to_signed(-46,32);
--			when -723 => sin_inv_data <= to_signed(-46,32);
--			when -722 => sin_inv_data <= to_signed(-46,32);
--			when -721 => sin_inv_data <= to_signed(-46,32);
--			when -720 => sin_inv_data <= to_signed(-46,32);
--			when -719 => sin_inv_data <= to_signed(-46,32);
--			when -718 => sin_inv_data <= to_signed(-46,32);
--			when -717 => sin_inv_data <= to_signed(-46,32);
--			when -716 => sin_inv_data <= to_signed(-46,32);
--			when -715 => sin_inv_data <= to_signed(-46,32);
--			when -714 => sin_inv_data <= to_signed(-46,32);
--			when -713 => sin_inv_data <= to_signed(-45,32);
--			when -712 => sin_inv_data <= to_signed(-45,32);
--			when -711 => sin_inv_data <= to_signed(-45,32);
--			when -710 => sin_inv_data <= to_signed(-45,32);
--			when -709 => sin_inv_data <= to_signed(-45,32);
--			when -708 => sin_inv_data <= to_signed(-45,32);
--			when -707 => sin_inv_data <= to_signed(-45,32);
--			when -706 => sin_inv_data <= to_signed(-45,32);
--			when -705 => sin_inv_data <= to_signed(-45,32);
--			when -704 => sin_inv_data <= to_signed(-45,32);
--			when -703 => sin_inv_data <= to_signed(-45,32);
--			when -702 => sin_inv_data <= to_signed(-45,32);
--			when -701 => sin_inv_data <= to_signed(-45,32);
--			when -700 => sin_inv_data <= to_signed(-44,32);
--			when -699 => sin_inv_data <= to_signed(-44,32);
--			when -698 => sin_inv_data <= to_signed(-44,32);
--			when -697 => sin_inv_data <= to_signed(-44,32);
--			when -696 => sin_inv_data <= to_signed(-44,32);
--			when -695 => sin_inv_data <= to_signed(-44,32);
--			when -694 => sin_inv_data <= to_signed(-44,32);
--			when -693 => sin_inv_data <= to_signed(-44,32);
--			when -692 => sin_inv_data <= to_signed(-44,32);
--			when -691 => sin_inv_data <= to_signed(-44,32);
--			when -690 => sin_inv_data <= to_signed(-44,32);
--			when -689 => sin_inv_data <= to_signed(-44,32);
--			when -688 => sin_inv_data <= to_signed(-43,32);
--			when -687 => sin_inv_data <= to_signed(-43,32);
--			when -686 => sin_inv_data <= to_signed(-43,32);
--			when -685 => sin_inv_data <= to_signed(-43,32);
--			when -684 => sin_inv_data <= to_signed(-43,32);
--			when -683 => sin_inv_data <= to_signed(-43,32);
--			when -682 => sin_inv_data <= to_signed(-43,32);
--			when -681 => sin_inv_data <= to_signed(-43,32);
--			when -680 => sin_inv_data <= to_signed(-43,32);
--			when -679 => sin_inv_data <= to_signed(-43,32);
--			when -678 => sin_inv_data <= to_signed(-43,32);
--			when -677 => sin_inv_data <= to_signed(-43,32);
--			when -676 => sin_inv_data <= to_signed(-43,32);
--			when -675 => sin_inv_data <= to_signed(-42,32);
--			when -674 => sin_inv_data <= to_signed(-42,32);
--			when -673 => sin_inv_data <= to_signed(-42,32);
--			when -672 => sin_inv_data <= to_signed(-42,32);
--			when -671 => sin_inv_data <= to_signed(-42,32);
--			when -670 => sin_inv_data <= to_signed(-42,32);
--			when -669 => sin_inv_data <= to_signed(-42,32);
--			when -668 => sin_inv_data <= to_signed(-42,32);
--			when -667 => sin_inv_data <= to_signed(-42,32);
--			when -666 => sin_inv_data <= to_signed(-42,32);
--			when -665 => sin_inv_data <= to_signed(-42,32);
--			when -664 => sin_inv_data <= to_signed(-42,32);
--			when -663 => sin_inv_data <= to_signed(-42,32);
--			when -662 => sin_inv_data <= to_signed(-41,32);
--			when -661 => sin_inv_data <= to_signed(-41,32);
--			when -660 => sin_inv_data <= to_signed(-41,32);
--			when -659 => sin_inv_data <= to_signed(-41,32);
--			when -658 => sin_inv_data <= to_signed(-41,32);
--			when -657 => sin_inv_data <= to_signed(-41,32);
--			when -656 => sin_inv_data <= to_signed(-41,32);
--			when -655 => sin_inv_data <= to_signed(-41,32);
--			when -654 => sin_inv_data <= to_signed(-41,32);
--			when -653 => sin_inv_data <= to_signed(-41,32);
--			when -652 => sin_inv_data <= to_signed(-41,32);
--			when -651 => sin_inv_data <= to_signed(-41,32);
--			when -650 => sin_inv_data <= to_signed(-41,32);
--			when -649 => sin_inv_data <= to_signed(-40,32);
--			when -648 => sin_inv_data <= to_signed(-40,32);
--			when -647 => sin_inv_data <= to_signed(-40,32);
--			when -646 => sin_inv_data <= to_signed(-40,32);
--			when -645 => sin_inv_data <= to_signed(-40,32);
--			when -644 => sin_inv_data <= to_signed(-40,32);
--			when -643 => sin_inv_data <= to_signed(-40,32);
--			when -642 => sin_inv_data <= to_signed(-40,32);
--			when -641 => sin_inv_data <= to_signed(-40,32);
--			when -640 => sin_inv_data <= to_signed(-40,32);
--			when -639 => sin_inv_data <= to_signed(-40,32);
--			when -638 => sin_inv_data <= to_signed(-40,32);
--			when -637 => sin_inv_data <= to_signed(-40,32);
--			when -636 => sin_inv_data <= to_signed(-39,32);
--			when -635 => sin_inv_data <= to_signed(-39,32);
--			when -634 => sin_inv_data <= to_signed(-39,32);
--			when -633 => sin_inv_data <= to_signed(-39,32);
--			when -632 => sin_inv_data <= to_signed(-39,32);
--			when -631 => sin_inv_data <= to_signed(-39,32);
--			when -630 => sin_inv_data <= to_signed(-39,32);
--			when -629 => sin_inv_data <= to_signed(-39,32);
--			when -628 => sin_inv_data <= to_signed(-39,32);
--			when -627 => sin_inv_data <= to_signed(-39,32);
--			when -626 => sin_inv_data <= to_signed(-39,32);
--			when -625 => sin_inv_data <= to_signed(-39,32);
--			when -624 => sin_inv_data <= to_signed(-39,32);
--			when -623 => sin_inv_data <= to_signed(-39,32);
--			when -622 => sin_inv_data <= to_signed(-38,32);
--			when -621 => sin_inv_data <= to_signed(-38,32);
--			when -620 => sin_inv_data <= to_signed(-38,32);
--			when -619 => sin_inv_data <= to_signed(-38,32);
--			when -618 => sin_inv_data <= to_signed(-38,32);
--			when -617 => sin_inv_data <= to_signed(-38,32);
--			when -616 => sin_inv_data <= to_signed(-38,32);
--			when -615 => sin_inv_data <= to_signed(-38,32);
--			when -614 => sin_inv_data <= to_signed(-38,32);
--			when -613 => sin_inv_data <= to_signed(-38,32);
--			when -612 => sin_inv_data <= to_signed(-38,32);
--			when -611 => sin_inv_data <= to_signed(-38,32);
--			when -610 => sin_inv_data <= to_signed(-38,32);
--			when -609 => sin_inv_data <= to_signed(-38,32);
--			when -608 => sin_inv_data <= to_signed(-37,32);
--			when -607 => sin_inv_data <= to_signed(-37,32);
--			when -606 => sin_inv_data <= to_signed(-37,32);
--			when -605 => sin_inv_data <= to_signed(-37,32);
--			when -604 => sin_inv_data <= to_signed(-37,32);
--			when -603 => sin_inv_data <= to_signed(-37,32);
--			when -602 => sin_inv_data <= to_signed(-37,32);
--			when -601 => sin_inv_data <= to_signed(-37,32);
--			when -600 => sin_inv_data <= to_signed(-37,32);
--			when -599 => sin_inv_data <= to_signed(-37,32);
--			when -598 => sin_inv_data <= to_signed(-37,32);
--			when -597 => sin_inv_data <= to_signed(-37,32);
--			when -596 => sin_inv_data <= to_signed(-37,32);
--			when -595 => sin_inv_data <= to_signed(-37,32);
--			when -594 => sin_inv_data <= to_signed(-36,32);
--			when -593 => sin_inv_data <= to_signed(-36,32);
--			when -592 => sin_inv_data <= to_signed(-36,32);
--			when -591 => sin_inv_data <= to_signed(-36,32);
--			when -590 => sin_inv_data <= to_signed(-36,32);
--			when -589 => sin_inv_data <= to_signed(-36,32);
--			when -588 => sin_inv_data <= to_signed(-36,32);
--			when -587 => sin_inv_data <= to_signed(-36,32);
--			when -586 => sin_inv_data <= to_signed(-36,32);
--			when -585 => sin_inv_data <= to_signed(-36,32);
--			when -584 => sin_inv_data <= to_signed(-36,32);
--			when -583 => sin_inv_data <= to_signed(-36,32);
--			when -582 => sin_inv_data <= to_signed(-36,32);
--			when -581 => sin_inv_data <= to_signed(-36,32);
--			when -580 => sin_inv_data <= to_signed(-35,32);
--			when -579 => sin_inv_data <= to_signed(-35,32);
--			when -578 => sin_inv_data <= to_signed(-35,32);
--			when -577 => sin_inv_data <= to_signed(-35,32);
--			when -576 => sin_inv_data <= to_signed(-35,32);
--			when -575 => sin_inv_data <= to_signed(-35,32);
--			when -574 => sin_inv_data <= to_signed(-35,32);
--			when -573 => sin_inv_data <= to_signed(-35,32);
--			when -572 => sin_inv_data <= to_signed(-35,32);
--			when -571 => sin_inv_data <= to_signed(-35,32);
--			when -570 => sin_inv_data <= to_signed(-35,32);
--			when -569 => sin_inv_data <= to_signed(-35,32);
--			when -568 => sin_inv_data <= to_signed(-35,32);
--			when -567 => sin_inv_data <= to_signed(-35,32);
--			when -566 => sin_inv_data <= to_signed(-34,32);
--			when -565 => sin_inv_data <= to_signed(-34,32);
--			when -564 => sin_inv_data <= to_signed(-34,32);
--			when -563 => sin_inv_data <= to_signed(-34,32);
--			when -562 => sin_inv_data <= to_signed(-34,32);
--			when -561 => sin_inv_data <= to_signed(-34,32);
--			when -560 => sin_inv_data <= to_signed(-34,32);
--			when -559 => sin_inv_data <= to_signed(-34,32);
--			when -558 => sin_inv_data <= to_signed(-34,32);
--			when -557 => sin_inv_data <= to_signed(-34,32);
--			when -556 => sin_inv_data <= to_signed(-34,32);
--			when -555 => sin_inv_data <= to_signed(-34,32);
--			when -554 => sin_inv_data <= to_signed(-34,32);
--			when -553 => sin_inv_data <= to_signed(-34,32);
--			when -552 => sin_inv_data <= to_signed(-34,32);
--			when -551 => sin_inv_data <= to_signed(-33,32);
--			when -550 => sin_inv_data <= to_signed(-33,32);
--			when -549 => sin_inv_data <= to_signed(-33,32);
--			when -548 => sin_inv_data <= to_signed(-33,32);
--			when -547 => sin_inv_data <= to_signed(-33,32);
--			when -546 => sin_inv_data <= to_signed(-33,32);
--			when -545 => sin_inv_data <= to_signed(-33,32);
--			when -544 => sin_inv_data <= to_signed(-33,32);
--			when -543 => sin_inv_data <= to_signed(-33,32);
--			when -542 => sin_inv_data <= to_signed(-33,32);
--			when -541 => sin_inv_data <= to_signed(-33,32);
--			when -540 => sin_inv_data <= to_signed(-33,32);
--			when -539 => sin_inv_data <= to_signed(-33,32);
--			when -538 => sin_inv_data <= to_signed(-33,32);
--			when -537 => sin_inv_data <= to_signed(-32,32);
--			when -536 => sin_inv_data <= to_signed(-32,32);
--			when -535 => sin_inv_data <= to_signed(-32,32);
--			when -534 => sin_inv_data <= to_signed(-32,32);
--			when -533 => sin_inv_data <= to_signed(-32,32);
--			when -532 => sin_inv_data <= to_signed(-32,32);
--			when -531 => sin_inv_data <= to_signed(-32,32);
--			when -530 => sin_inv_data <= to_signed(-32,32);
--			when -529 => sin_inv_data <= to_signed(-32,32);
--			when -528 => sin_inv_data <= to_signed(-32,32);
--			when -527 => sin_inv_data <= to_signed(-32,32);
--			when -526 => sin_inv_data <= to_signed(-32,32);
--			when -525 => sin_inv_data <= to_signed(-32,32);
--			when -524 => sin_inv_data <= to_signed(-32,32);
--			when -523 => sin_inv_data <= to_signed(-32,32);
--			when -522 => sin_inv_data <= to_signed(-31,32);
--			when -521 => sin_inv_data <= to_signed(-31,32);
--			when -520 => sin_inv_data <= to_signed(-31,32);
--			when -519 => sin_inv_data <= to_signed(-31,32);
--			when -518 => sin_inv_data <= to_signed(-31,32);
--			when -517 => sin_inv_data <= to_signed(-31,32);
--			when -516 => sin_inv_data <= to_signed(-31,32);
--			when -515 => sin_inv_data <= to_signed(-31,32);
--			when -514 => sin_inv_data <= to_signed(-31,32);
--			when -513 => sin_inv_data <= to_signed(-31,32);
--			when -512 => sin_inv_data <= to_signed(-31,32);
--			when -511 => sin_inv_data <= to_signed(-31,32);
--			when -510 => sin_inv_data <= to_signed(-31,32);
--			when -509 => sin_inv_data <= to_signed(-31,32);
--			when -508 => sin_inv_data <= to_signed(-31,32);
--			when -507 => sin_inv_data <= to_signed(-30,32);
--			when -506 => sin_inv_data <= to_signed(-30,32);
--			when -505 => sin_inv_data <= to_signed(-30,32);
--			when -504 => sin_inv_data <= to_signed(-30,32);
--			when -503 => sin_inv_data <= to_signed(-30,32);
--			when -502 => sin_inv_data <= to_signed(-30,32);
--			when -501 => sin_inv_data <= to_signed(-30,32);
--			when -500 => sin_inv_data <= to_signed(-30,32);
--			when -499 => sin_inv_data <= to_signed(-30,32);
--			when -498 => sin_inv_data <= to_signed(-30,32);
--			when -497 => sin_inv_data <= to_signed(-30,32);
--			when -496 => sin_inv_data <= to_signed(-30,32);
--			when -495 => sin_inv_data <= to_signed(-30,32);
--			when -494 => sin_inv_data <= to_signed(-30,32);
--			when -493 => sin_inv_data <= to_signed(-30,32);
--			when -492 => sin_inv_data <= to_signed(-29,32);
--			when -491 => sin_inv_data <= to_signed(-29,32);
--			when -490 => sin_inv_data <= to_signed(-29,32);
--			when -489 => sin_inv_data <= to_signed(-29,32);
--			when -488 => sin_inv_data <= to_signed(-29,32);
--			when -487 => sin_inv_data <= to_signed(-29,32);
--			when -486 => sin_inv_data <= to_signed(-29,32);
--			when -485 => sin_inv_data <= to_signed(-29,32);
--			when -484 => sin_inv_data <= to_signed(-29,32);
--			when -483 => sin_inv_data <= to_signed(-29,32);
--			when -482 => sin_inv_data <= to_signed(-29,32);
--			when -481 => sin_inv_data <= to_signed(-29,32);
--			when -480 => sin_inv_data <= to_signed(-29,32);
--			when -479 => sin_inv_data <= to_signed(-29,32);
--			when -478 => sin_inv_data <= to_signed(-29,32);
--			when -477 => sin_inv_data <= to_signed(-28,32);
--			when -476 => sin_inv_data <= to_signed(-28,32);
--			when -475 => sin_inv_data <= to_signed(-28,32);
--			when -474 => sin_inv_data <= to_signed(-28,32);
--			when -473 => sin_inv_data <= to_signed(-28,32);
--			when -472 => sin_inv_data <= to_signed(-28,32);
--			when -471 => sin_inv_data <= to_signed(-28,32);
--			when -470 => sin_inv_data <= to_signed(-28,32);
--			when -469 => sin_inv_data <= to_signed(-28,32);
--			when -468 => sin_inv_data <= to_signed(-28,32);
--			when -467 => sin_inv_data <= to_signed(-28,32);
--			when -466 => sin_inv_data <= to_signed(-28,32);
--			when -465 => sin_inv_data <= to_signed(-28,32);
--			when -464 => sin_inv_data <= to_signed(-28,32);
--			when -463 => sin_inv_data <= to_signed(-28,32);
--			when -462 => sin_inv_data <= to_signed(-28,32);
--			when -461 => sin_inv_data <= to_signed(-27,32);
--			when -460 => sin_inv_data <= to_signed(-27,32);
--			when -459 => sin_inv_data <= to_signed(-27,32);
--			when -458 => sin_inv_data <= to_signed(-27,32);
--			when -457 => sin_inv_data <= to_signed(-27,32);
--			when -456 => sin_inv_data <= to_signed(-27,32);
--			when -455 => sin_inv_data <= to_signed(-27,32);
--			when -454 => sin_inv_data <= to_signed(-27,32);
--			when -453 => sin_inv_data <= to_signed(-27,32);
--			when -452 => sin_inv_data <= to_signed(-27,32);
--			when -451 => sin_inv_data <= to_signed(-27,32);
--			when -450 => sin_inv_data <= to_signed(-27,32);
--			when -449 => sin_inv_data <= to_signed(-27,32);
--			when -448 => sin_inv_data <= to_signed(-27,32);
--			when -447 => sin_inv_data <= to_signed(-27,32);
--			when -446 => sin_inv_data <= to_signed(-26,32);
--			when -445 => sin_inv_data <= to_signed(-26,32);
--			when -444 => sin_inv_data <= to_signed(-26,32);
--			when -443 => sin_inv_data <= to_signed(-26,32);
--			when -442 => sin_inv_data <= to_signed(-26,32);
--			when -441 => sin_inv_data <= to_signed(-26,32);
--			when -440 => sin_inv_data <= to_signed(-26,32);
--			when -439 => sin_inv_data <= to_signed(-26,32);
--			when -438 => sin_inv_data <= to_signed(-26,32);
--			when -437 => sin_inv_data <= to_signed(-26,32);
--			when -436 => sin_inv_data <= to_signed(-26,32);
--			when -435 => sin_inv_data <= to_signed(-26,32);
--			when -434 => sin_inv_data <= to_signed(-26,32);
--			when -433 => sin_inv_data <= to_signed(-26,32);
--			when -432 => sin_inv_data <= to_signed(-26,32);
--			when -431 => sin_inv_data <= to_signed(-26,32);
--			when -430 => sin_inv_data <= to_signed(-25,32);
--			when -429 => sin_inv_data <= to_signed(-25,32);
--			when -428 => sin_inv_data <= to_signed(-25,32);
--			when -427 => sin_inv_data <= to_signed(-25,32);
--			when -426 => sin_inv_data <= to_signed(-25,32);
--			when -425 => sin_inv_data <= to_signed(-25,32);
--			when -424 => sin_inv_data <= to_signed(-25,32);
--			when -423 => sin_inv_data <= to_signed(-25,32);
--			when -422 => sin_inv_data <= to_signed(-25,32);
--			when -421 => sin_inv_data <= to_signed(-25,32);
--			when -420 => sin_inv_data <= to_signed(-25,32);
--			when -419 => sin_inv_data <= to_signed(-25,32);
--			when -418 => sin_inv_data <= to_signed(-25,32);
--			when -417 => sin_inv_data <= to_signed(-25,32);
--			when -416 => sin_inv_data <= to_signed(-25,32);
--			when -415 => sin_inv_data <= to_signed(-25,32);
--			when -414 => sin_inv_data <= to_signed(-24,32);
--			when -413 => sin_inv_data <= to_signed(-24,32);
--			when -412 => sin_inv_data <= to_signed(-24,32);
--			when -411 => sin_inv_data <= to_signed(-24,32);
--			when -410 => sin_inv_data <= to_signed(-24,32);
--			when -409 => sin_inv_data <= to_signed(-24,32);
--			when -408 => sin_inv_data <= to_signed(-24,32);
--			when -407 => sin_inv_data <= to_signed(-24,32);
--			when -406 => sin_inv_data <= to_signed(-24,32);
--			when -405 => sin_inv_data <= to_signed(-24,32);
--			when -404 => sin_inv_data <= to_signed(-24,32);
--			when -403 => sin_inv_data <= to_signed(-24,32);
--			when -402 => sin_inv_data <= to_signed(-24,32);
--			when -401 => sin_inv_data <= to_signed(-24,32);
--			when -400 => sin_inv_data <= to_signed(-24,32);
--			when -399 => sin_inv_data <= to_signed(-24,32);
--			when -398 => sin_inv_data <= to_signed(-23,32);
--			when -397 => sin_inv_data <= to_signed(-23,32);
--			when -396 => sin_inv_data <= to_signed(-23,32);
--			when -395 => sin_inv_data <= to_signed(-23,32);
--			when -394 => sin_inv_data <= to_signed(-23,32);
--			when -393 => sin_inv_data <= to_signed(-23,32);
--			when -392 => sin_inv_data <= to_signed(-23,32);
--			when -391 => sin_inv_data <= to_signed(-23,32);
--			when -390 => sin_inv_data <= to_signed(-23,32);
--			when -389 => sin_inv_data <= to_signed(-23,32);
--			when -388 => sin_inv_data <= to_signed(-23,32);
--			when -387 => sin_inv_data <= to_signed(-23,32);
--			when -386 => sin_inv_data <= to_signed(-23,32);
--			when -385 => sin_inv_data <= to_signed(-23,32);
--			when -384 => sin_inv_data <= to_signed(-23,32);
--			when -383 => sin_inv_data <= to_signed(-23,32);
--			when -382 => sin_inv_data <= to_signed(-22,32);
--			when -381 => sin_inv_data <= to_signed(-22,32);
--			when -380 => sin_inv_data <= to_signed(-22,32);
--			when -379 => sin_inv_data <= to_signed(-22,32);
--			when -378 => sin_inv_data <= to_signed(-22,32);
--			when -377 => sin_inv_data <= to_signed(-22,32);
--			when -376 => sin_inv_data <= to_signed(-22,32);
--			when -375 => sin_inv_data <= to_signed(-22,32);
--			when -374 => sin_inv_data <= to_signed(-22,32);
--			when -373 => sin_inv_data <= to_signed(-22,32);
--			when -372 => sin_inv_data <= to_signed(-22,32);
--			when -371 => sin_inv_data <= to_signed(-22,32);
--			when -370 => sin_inv_data <= to_signed(-22,32);
--			when -369 => sin_inv_data <= to_signed(-22,32);
--			when -368 => sin_inv_data <= to_signed(-22,32);
--			when -367 => sin_inv_data <= to_signed(-22,32);
--			when -366 => sin_inv_data <= to_signed(-21,32);
--			when -365 => sin_inv_data <= to_signed(-21,32);
--			when -364 => sin_inv_data <= to_signed(-21,32);
--			when -363 => sin_inv_data <= to_signed(-21,32);
--			when -362 => sin_inv_data <= to_signed(-21,32);
--			when -361 => sin_inv_data <= to_signed(-21,32);
--			when -360 => sin_inv_data <= to_signed(-21,32);
--			when -359 => sin_inv_data <= to_signed(-21,32);
--			when -358 => sin_inv_data <= to_signed(-21,32);
--			when -357 => sin_inv_data <= to_signed(-21,32);
--			when -356 => sin_inv_data <= to_signed(-21,32);
--			when -355 => sin_inv_data <= to_signed(-21,32);
--			when -354 => sin_inv_data <= to_signed(-21,32);
--			when -353 => sin_inv_data <= to_signed(-21,32);
--			when -352 => sin_inv_data <= to_signed(-21,32);
--			when -351 => sin_inv_data <= to_signed(-21,32);
--			when -350 => sin_inv_data <= to_signed(-20,32);
--			when -349 => sin_inv_data <= to_signed(-20,32);
--			when -348 => sin_inv_data <= to_signed(-20,32);
--			when -347 => sin_inv_data <= to_signed(-20,32);
--			when -346 => sin_inv_data <= to_signed(-20,32);
--			when -345 => sin_inv_data <= to_signed(-20,32);
--			when -344 => sin_inv_data <= to_signed(-20,32);
--			when -343 => sin_inv_data <= to_signed(-20,32);
--			when -342 => sin_inv_data <= to_signed(-20,32);
--			when -341 => sin_inv_data <= to_signed(-20,32);
--			when -340 => sin_inv_data <= to_signed(-20,32);
--			when -339 => sin_inv_data <= to_signed(-20,32);
--			when -338 => sin_inv_data <= to_signed(-20,32);
--			when -337 => sin_inv_data <= to_signed(-20,32);
--			when -336 => sin_inv_data <= to_signed(-20,32);
--			when -335 => sin_inv_data <= to_signed(-20,32);
--			when -334 => sin_inv_data <= to_signed(-20,32);
--			when -333 => sin_inv_data <= to_signed(-19,32);
--			when -332 => sin_inv_data <= to_signed(-19,32);
--			when -331 => sin_inv_data <= to_signed(-19,32);
--			when -330 => sin_inv_data <= to_signed(-19,32);
--			when -329 => sin_inv_data <= to_signed(-19,32);
--			when -328 => sin_inv_data <= to_signed(-19,32);
--			when -327 => sin_inv_data <= to_signed(-19,32);
--			when -326 => sin_inv_data <= to_signed(-19,32);
--			when -325 => sin_inv_data <= to_signed(-19,32);
--			when -324 => sin_inv_data <= to_signed(-19,32);
--			when -323 => sin_inv_data <= to_signed(-19,32);
--			when -322 => sin_inv_data <= to_signed(-19,32);
--			when -321 => sin_inv_data <= to_signed(-19,32);
--			when -320 => sin_inv_data <= to_signed(-19,32);
--			when -319 => sin_inv_data <= to_signed(-19,32);
--			when -318 => sin_inv_data <= to_signed(-19,32);
--			when -317 => sin_inv_data <= to_signed(-18,32);
--			when -316 => sin_inv_data <= to_signed(-18,32);
--			when -315 => sin_inv_data <= to_signed(-18,32);
--			when -314 => sin_inv_data <= to_signed(-18,32);
--			when -313 => sin_inv_data <= to_signed(-18,32);
--			when -312 => sin_inv_data <= to_signed(-18,32);
--			when -311 => sin_inv_data <= to_signed(-18,32);
--			when -310 => sin_inv_data <= to_signed(-18,32);
--			when -309 => sin_inv_data <= to_signed(-18,32);
--			when -308 => sin_inv_data <= to_signed(-18,32);
--			when -307 => sin_inv_data <= to_signed(-18,32);
--			when -306 => sin_inv_data <= to_signed(-18,32);
--			when -305 => sin_inv_data <= to_signed(-18,32);
--			when -304 => sin_inv_data <= to_signed(-18,32);
--			when -303 => sin_inv_data <= to_signed(-18,32);
--			when -302 => sin_inv_data <= to_signed(-18,32);
--			when -301 => sin_inv_data <= to_signed(-18,32);
--			when -300 => sin_inv_data <= to_signed(-17,32);
--			when -299 => sin_inv_data <= to_signed(-17,32);
--			when -298 => sin_inv_data <= to_signed(-17,32);
--			when -297 => sin_inv_data <= to_signed(-17,32);
--			when -296 => sin_inv_data <= to_signed(-17,32);
--			when -295 => sin_inv_data <= to_signed(-17,32);
--			when -294 => sin_inv_data <= to_signed(-17,32);
--			when -293 => sin_inv_data <= to_signed(-17,32);
--			when -292 => sin_inv_data <= to_signed(-17,32);
--			when -291 => sin_inv_data <= to_signed(-17,32);
--			when -290 => sin_inv_data <= to_signed(-17,32);
--			when -289 => sin_inv_data <= to_signed(-17,32);
--			when -288 => sin_inv_data <= to_signed(-17,32);
--			when -287 => sin_inv_data <= to_signed(-17,32);
--			when -286 => sin_inv_data <= to_signed(-17,32);
--			when -285 => sin_inv_data <= to_signed(-17,32);
--			when -284 => sin_inv_data <= to_signed(-16,32);
--			when -283 => sin_inv_data <= to_signed(-16,32);
--			when -282 => sin_inv_data <= to_signed(-16,32);
--			when -281 => sin_inv_data <= to_signed(-16,32);
--			when -280 => sin_inv_data <= to_signed(-16,32);
--			when -279 => sin_inv_data <= to_signed(-16,32);
--			when -278 => sin_inv_data <= to_signed(-16,32);
--			when -277 => sin_inv_data <= to_signed(-16,32);
--			when -276 => sin_inv_data <= to_signed(-16,32);
--			when -275 => sin_inv_data <= to_signed(-16,32);
--			when -274 => sin_inv_data <= to_signed(-16,32);
--			when -273 => sin_inv_data <= to_signed(-16,32);
--			when -272 => sin_inv_data <= to_signed(-16,32);
--			when -271 => sin_inv_data <= to_signed(-16,32);
--			when -270 => sin_inv_data <= to_signed(-16,32);
--			when -269 => sin_inv_data <= to_signed(-16,32);
--			when -268 => sin_inv_data <= to_signed(-16,32);
--			when -267 => sin_inv_data <= to_signed(-15,32);
--			when -266 => sin_inv_data <= to_signed(-15,32);
--			when -265 => sin_inv_data <= to_signed(-15,32);
--			when -264 => sin_inv_data <= to_signed(-15,32);
--			when -263 => sin_inv_data <= to_signed(-15,32);
--			when -262 => sin_inv_data <= to_signed(-15,32);
--			when -261 => sin_inv_data <= to_signed(-15,32);
--			when -260 => sin_inv_data <= to_signed(-15,32);
--			when -259 => sin_inv_data <= to_signed(-15,32);
--			when -258 => sin_inv_data <= to_signed(-15,32);
--			when -257 => sin_inv_data <= to_signed(-15,32);
--			when -256 => sin_inv_data <= to_signed(-15,32);
--			when -255 => sin_inv_data <= to_signed(-15,32);
--			when -254 => sin_inv_data <= to_signed(-15,32);
--			when -253 => sin_inv_data <= to_signed(-15,32);
--			when -252 => sin_inv_data <= to_signed(-15,32);
--			when -251 => sin_inv_data <= to_signed(-15,32);
--			when -250 => sin_inv_data <= to_signed(-14,32);
--			when -249 => sin_inv_data <= to_signed(-14,32);
--			when -248 => sin_inv_data <= to_signed(-14,32);
--			when -247 => sin_inv_data <= to_signed(-14,32);
--			when -246 => sin_inv_data <= to_signed(-14,32);
--			when -245 => sin_inv_data <= to_signed(-14,32);
--			when -244 => sin_inv_data <= to_signed(-14,32);
--			when -243 => sin_inv_data <= to_signed(-14,32);
--			when -242 => sin_inv_data <= to_signed(-14,32);
--			when -241 => sin_inv_data <= to_signed(-14,32);
--			when -240 => sin_inv_data <= to_signed(-14,32);
--			when -239 => sin_inv_data <= to_signed(-14,32);
--			when -238 => sin_inv_data <= to_signed(-14,32);
--			when -237 => sin_inv_data <= to_signed(-14,32);
--			when -236 => sin_inv_data <= to_signed(-14,32);
--			when -235 => sin_inv_data <= to_signed(-14,32);
--			when -234 => sin_inv_data <= to_signed(-14,32);
--			when -233 => sin_inv_data <= to_signed(-13,32);
--			when -232 => sin_inv_data <= to_signed(-13,32);
--			when -231 => sin_inv_data <= to_signed(-13,32);
--			when -230 => sin_inv_data <= to_signed(-13,32);
--			when -229 => sin_inv_data <= to_signed(-13,32);
--			when -228 => sin_inv_data <= to_signed(-13,32);
--			when -227 => sin_inv_data <= to_signed(-13,32);
--			when -226 => sin_inv_data <= to_signed(-13,32);
--			when -225 => sin_inv_data <= to_signed(-13,32);
--			when -224 => sin_inv_data <= to_signed(-13,32);
--			when -223 => sin_inv_data <= to_signed(-13,32);
--			when -222 => sin_inv_data <= to_signed(-13,32);
--			when -221 => sin_inv_data <= to_signed(-13,32);
--			when -220 => sin_inv_data <= to_signed(-13,32);
--			when -219 => sin_inv_data <= to_signed(-13,32);
--			when -218 => sin_inv_data <= to_signed(-13,32);
--			when -217 => sin_inv_data <= to_signed(-13,32);
--			when -216 => sin_inv_data <= to_signed(-12,32);
--			when -215 => sin_inv_data <= to_signed(-12,32);
--			when -214 => sin_inv_data <= to_signed(-12,32);
--			when -213 => sin_inv_data <= to_signed(-12,32);
--			when -212 => sin_inv_data <= to_signed(-12,32);
--			when -211 => sin_inv_data <= to_signed(-12,32);
--			when -210 => sin_inv_data <= to_signed(-12,32);
--			when -209 => sin_inv_data <= to_signed(-12,32);
--			when -208 => sin_inv_data <= to_signed(-12,32);
--			when -207 => sin_inv_data <= to_signed(-12,32);
--			when -206 => sin_inv_data <= to_signed(-12,32);
--			when -205 => sin_inv_data <= to_signed(-12,32);
--			when -204 => sin_inv_data <= to_signed(-12,32);
--			when -203 => sin_inv_data <= to_signed(-12,32);
--			when -202 => sin_inv_data <= to_signed(-12,32);
--			when -201 => sin_inv_data <= to_signed(-12,32);
--			when -200 => sin_inv_data <= to_signed(-12,32);
--			when -199 => sin_inv_data <= to_signed(-11,32);
--			when -198 => sin_inv_data <= to_signed(-11,32);
--			when -197 => sin_inv_data <= to_signed(-11,32);
--			when -196 => sin_inv_data <= to_signed(-11,32);
--			when -195 => sin_inv_data <= to_signed(-11,32);
--			when -194 => sin_inv_data <= to_signed(-11,32);
--			when -193 => sin_inv_data <= to_signed(-11,32);
--			when -192 => sin_inv_data <= to_signed(-11,32);
--			when -191 => sin_inv_data <= to_signed(-11,32);
--			when -190 => sin_inv_data <= to_signed(-11,32);
--			when -189 => sin_inv_data <= to_signed(-11,32);
--			when -188 => sin_inv_data <= to_signed(-11,32);
--			when -187 => sin_inv_data <= to_signed(-11,32);
--			when -186 => sin_inv_data <= to_signed(-11,32);
--			when -185 => sin_inv_data <= to_signed(-11,32);
--			when -184 => sin_inv_data <= to_signed(-11,32);
--			when -183 => sin_inv_data <= to_signed(-11,32);
--			when -182 => sin_inv_data <= to_signed(-10,32);
--			when -181 => sin_inv_data <= to_signed(-10,32);
--			when -180 => sin_inv_data <= to_signed(-10,32);
--			when -179 => sin_inv_data <= to_signed(-10,32);
--			when -178 => sin_inv_data <= to_signed(-10,32);
--			when -177 => sin_inv_data <= to_signed(-10,32);
--			when -176 => sin_inv_data <= to_signed(-10,32);
--			when -175 => sin_inv_data <= to_signed(-10,32);
--			when -174 => sin_inv_data <= to_signed(-10,32);
--			when -173 => sin_inv_data <= to_signed(-10,32);
--			when -172 => sin_inv_data <= to_signed(-10,32);
--			when -171 => sin_inv_data <= to_signed(-10,32);
--			when -170 => sin_inv_data <= to_signed(-10,32);
--			when -169 => sin_inv_data <= to_signed(-10,32);
--			when -168 => sin_inv_data <= to_signed(-10,32);
--			when -167 => sin_inv_data <= to_signed(-10,32);
--			when -166 => sin_inv_data <= to_signed(-10,32);
--			when -165 => sin_inv_data <= to_signed(-9,32);
--			when -164 => sin_inv_data <= to_signed(-9,32);
--			when -163 => sin_inv_data <= to_signed(-9,32);
--			when -162 => sin_inv_data <= to_signed(-9,32);
--			when -161 => sin_inv_data <= to_signed(-9,32);
--			when -160 => sin_inv_data <= to_signed(-9,32);
--			when -159 => sin_inv_data <= to_signed(-9,32);
--			when -158 => sin_inv_data <= to_signed(-9,32);
--			when -157 => sin_inv_data <= to_signed(-9,32);
--			when -156 => sin_inv_data <= to_signed(-9,32);
--			when -155 => sin_inv_data <= to_signed(-9,32);
--			when -154 => sin_inv_data <= to_signed(-9,32);
--			when -153 => sin_inv_data <= to_signed(-9,32);
--			when -152 => sin_inv_data <= to_signed(-9,32);
--			when -151 => sin_inv_data <= to_signed(-9,32);
--			when -150 => sin_inv_data <= to_signed(-9,32);
--			when -149 => sin_inv_data <= to_signed(-9,32);
--			when -148 => sin_inv_data <= to_signed(-9,32);
--			when -147 => sin_inv_data <= to_signed(-8,32);
--			when -146 => sin_inv_data <= to_signed(-8,32);
--			when -145 => sin_inv_data <= to_signed(-8,32);
--			when -144 => sin_inv_data <= to_signed(-8,32);
--			when -143 => sin_inv_data <= to_signed(-8,32);
--			when -142 => sin_inv_data <= to_signed(-8,32);
--			when -141 => sin_inv_data <= to_signed(-8,32);
--			when -140 => sin_inv_data <= to_signed(-8,32);
--			when -139 => sin_inv_data <= to_signed(-8,32);
--			when -138 => sin_inv_data <= to_signed(-8,32);
--			when -137 => sin_inv_data <= to_signed(-8,32);
--			when -136 => sin_inv_data <= to_signed(-8,32);
--			when -135 => sin_inv_data <= to_signed(-8,32);
--			when -134 => sin_inv_data <= to_signed(-8,32);
--			when -133 => sin_inv_data <= to_signed(-8,32);
--			when -132 => sin_inv_data <= to_signed(-8,32);
--			when -131 => sin_inv_data <= to_signed(-8,32);
--			when -130 => sin_inv_data <= to_signed(-7,32);
--			when -129 => sin_inv_data <= to_signed(-7,32);
--			when -128 => sin_inv_data <= to_signed(-7,32);
--			when -127 => sin_inv_data <= to_signed(-7,32);
--			when -126 => sin_inv_data <= to_signed(-7,32);
--			when -125 => sin_inv_data <= to_signed(-7,32);
--			when -124 => sin_inv_data <= to_signed(-7,32);
--			when -123 => sin_inv_data <= to_signed(-7,32);
--			when -122 => sin_inv_data <= to_signed(-7,32);
--			when -121 => sin_inv_data <= to_signed(-7,32);
--			when -120 => sin_inv_data <= to_signed(-7,32);
--			when -119 => sin_inv_data <= to_signed(-7,32);
--			when -118 => sin_inv_data <= to_signed(-7,32);
--			when -117 => sin_inv_data <= to_signed(-7,32);
--			when -116 => sin_inv_data <= to_signed(-7,32);
--			when -115 => sin_inv_data <= to_signed(-7,32);
--			when -114 => sin_inv_data <= to_signed(-7,32);
--			when -113 => sin_inv_data <= to_signed(-6,32);
--			when -112 => sin_inv_data <= to_signed(-6,32);
--			when -111 => sin_inv_data <= to_signed(-6,32);
--			when -110 => sin_inv_data <= to_signed(-6,32);
--			when -109 => sin_inv_data <= to_signed(-6,32);
--			when -108 => sin_inv_data <= to_signed(-6,32);
--			when -107 => sin_inv_data <= to_signed(-6,32);
--			when -106 => sin_inv_data <= to_signed(-6,32);
--			when -105 => sin_inv_data <= to_signed(-6,32);
--			when -104 => sin_inv_data <= to_signed(-6,32);
--			when -103 => sin_inv_data <= to_signed(-6,32);
--			when -102 => sin_inv_data <= to_signed(-6,32);
--			when -101 => sin_inv_data <= to_signed(-6,32);
--			when -100 => sin_inv_data <= to_signed(-6,32);
--			when -99 => sin_inv_data <= to_signed(-6,32);
--			when -98 => sin_inv_data <= to_signed(-6,32);
--			when -97 => sin_inv_data <= to_signed(-6,32);
--			when -96 => sin_inv_data <= to_signed(-6,32);
--			when -95 => sin_inv_data <= to_signed(-5,32);
--			when -94 => sin_inv_data <= to_signed(-5,32);
--			when -93 => sin_inv_data <= to_signed(-5,32);
--			when -92 => sin_inv_data <= to_signed(-5,32);
--			when -91 => sin_inv_data <= to_signed(-5,32);
--			when -90 => sin_inv_data <= to_signed(-5,32);
--			when -89 => sin_inv_data <= to_signed(-5,32);
--			when -88 => sin_inv_data <= to_signed(-5,32);
--			when -87 => sin_inv_data <= to_signed(-5,32);
--			when -86 => sin_inv_data <= to_signed(-5,32);
--			when -85 => sin_inv_data <= to_signed(-5,32);
--			when -84 => sin_inv_data <= to_signed(-5,32);
--			when -83 => sin_inv_data <= to_signed(-5,32);
--			when -82 => sin_inv_data <= to_signed(-5,32);
--			when -81 => sin_inv_data <= to_signed(-5,32);
--			when -80 => sin_inv_data <= to_signed(-5,32);
--			when -79 => sin_inv_data <= to_signed(-5,32);
--			when -78 => sin_inv_data <= to_signed(-4,32);
--			when -77 => sin_inv_data <= to_signed(-4,32);
--			when -76 => sin_inv_data <= to_signed(-4,32);
--			when -75 => sin_inv_data <= to_signed(-4,32);
--			when -74 => sin_inv_data <= to_signed(-4,32);
--			when -73 => sin_inv_data <= to_signed(-4,32);
--			when -72 => sin_inv_data <= to_signed(-4,32);
--			when -71 => sin_inv_data <= to_signed(-4,32);
--			when -70 => sin_inv_data <= to_signed(-4,32);
--			when -69 => sin_inv_data <= to_signed(-4,32);
--			when -68 => sin_inv_data <= to_signed(-4,32);
--			when -67 => sin_inv_data <= to_signed(-4,32);
--			when -66 => sin_inv_data <= to_signed(-4,32);
--			when -65 => sin_inv_data <= to_signed(-4,32);
--			when -64 => sin_inv_data <= to_signed(-4,32);
--			when -63 => sin_inv_data <= to_signed(-4,32);
--			when -62 => sin_inv_data <= to_signed(-4,32);
--			when -61 => sin_inv_data <= to_signed(-3,32);
--			when -60 => sin_inv_data <= to_signed(-3,32);
--			when -59 => sin_inv_data <= to_signed(-3,32);
--			when -58 => sin_inv_data <= to_signed(-3,32);
--			when -57 => sin_inv_data <= to_signed(-3,32);
--			when -56 => sin_inv_data <= to_signed(-3,32);
--			when -55 => sin_inv_data <= to_signed(-3,32);
--			when -54 => sin_inv_data <= to_signed(-3,32);
--			when -53 => sin_inv_data <= to_signed(-3,32);
--			when -52 => sin_inv_data <= to_signed(-3,32);
--			when -51 => sin_inv_data <= to_signed(-3,32);
--			when -50 => sin_inv_data <= to_signed(-3,32);
--			when -49 => sin_inv_data <= to_signed(-3,32);
--			when -48 => sin_inv_data <= to_signed(-3,32);
--			when -47 => sin_inv_data <= to_signed(-3,32);
--			when -46 => sin_inv_data <= to_signed(-3,32);
--			when -45 => sin_inv_data <= to_signed(-3,32);
--			when -44 => sin_inv_data <= to_signed(-3,32);
--			when -43 => sin_inv_data <= to_signed(-2,32);
--			when -42 => sin_inv_data <= to_signed(-2,32);
--			when -41 => sin_inv_data <= to_signed(-2,32);
--			when -40 => sin_inv_data <= to_signed(-2,32);
--			when -39 => sin_inv_data <= to_signed(-2,32);
--			when -38 => sin_inv_data <= to_signed(-2,32);
--			when -37 => sin_inv_data <= to_signed(-2,32);
--			when -36 => sin_inv_data <= to_signed(-2,32);
--			when -35 => sin_inv_data <= to_signed(-2,32);
--			when -34 => sin_inv_data <= to_signed(-2,32);
--			when -33 => sin_inv_data <= to_signed(-2,32);
--			when -32 => sin_inv_data <= to_signed(-2,32);
--			when -31 => sin_inv_data <= to_signed(-2,32);
--			when -30 => sin_inv_data <= to_signed(-2,32);
--			when -29 => sin_inv_data <= to_signed(-2,32);
--			when -28 => sin_inv_data <= to_signed(-2,32);
--			when -27 => sin_inv_data <= to_signed(-2,32);
--			when -26 => sin_inv_data <= to_signed(-1,32);
--			when -25 => sin_inv_data <= to_signed(-1,32);
--			when -24 => sin_inv_data <= to_signed(-1,32);
--			when -23 => sin_inv_data <= to_signed(-1,32);
--			when -22 => sin_inv_data <= to_signed(-1,32);
--			when -21 => sin_inv_data <= to_signed(-1,32);
--			when -20 => sin_inv_data <= to_signed(-1,32);
--			when -19 => sin_inv_data <= to_signed(-1,32);
--			when -18 => sin_inv_data <= to_signed(-1,32);
--			when -17 => sin_inv_data <= to_signed(-1,32);
--			when -16 => sin_inv_data <= to_signed(-1,32);
--			when -15 => sin_inv_data <= to_signed(-1,32);
--			when -14 => sin_inv_data <= to_signed(-1,32);
--			when -13 => sin_inv_data <= to_signed(-1,32);
--			when -12 => sin_inv_data <= to_signed(-1,32);
--			when -11 => sin_inv_data <= to_signed(-1,32);
--			when -10 => sin_inv_data <= to_signed(-1,32);
--			when -9 => sin_inv_data <= to_signed(-1,32);
--			when -8 => sin_inv_data <= to_signed(0,32);
--			when -7 => sin_inv_data <= to_signed(0,32);
--			when -6 => sin_inv_data <= to_signed(0,32);
--			when -5 => sin_inv_data <= to_signed(0,32);
--			when -4 => sin_inv_data <= to_signed(0,32);
--			when -3 => sin_inv_data <= to_signed(0,32);
--			when -2 => sin_inv_data <= to_signed(0,32);
--			when -1 => sin_inv_data <= to_signed(0,32);
--			when 0 => sin_inv_data <= to_signed(0,32);
--			when 1 => sin_inv_data <= to_signed(0,32);
--			when 2 => sin_inv_data <= to_signed(0,32);
--			when 3 => sin_inv_data <= to_signed(0,32);
--			when 4 => sin_inv_data <= to_signed(0,32);
--			when 5 => sin_inv_data <= to_signed(0,32);
--			when 6 => sin_inv_data <= to_signed(0,32);
--			when 7 => sin_inv_data <= to_signed(0,32);
--			when 8 => sin_inv_data <= to_signed(0,32);
--			when 9 => sin_inv_data <= to_signed(1,32);
--			when 10 => sin_inv_data <= to_signed(1,32);
--			when 11 => sin_inv_data <= to_signed(1,32);
--			when 12 => sin_inv_data <= to_signed(1,32);
--			when 13 => sin_inv_data <= to_signed(1,32);
--			when 14 => sin_inv_data <= to_signed(1,32);
--			when 15 => sin_inv_data <= to_signed(1,32);
--			when 16 => sin_inv_data <= to_signed(1,32);
--			when 17 => sin_inv_data <= to_signed(1,32);
--			when 18 => sin_inv_data <= to_signed(1,32);
--			when 19 => sin_inv_data <= to_signed(1,32);
--			when 20 => sin_inv_data <= to_signed(1,32);
--			when 21 => sin_inv_data <= to_signed(1,32);
--			when 22 => sin_inv_data <= to_signed(1,32);
--			when 23 => sin_inv_data <= to_signed(1,32);
--			when 24 => sin_inv_data <= to_signed(1,32);
--			when 25 => sin_inv_data <= to_signed(1,32);
--			when 26 => sin_inv_data <= to_signed(1,32);
--			when 27 => sin_inv_data <= to_signed(2,32);
--			when 28 => sin_inv_data <= to_signed(2,32);
--			when 29 => sin_inv_data <= to_signed(2,32);
--			when 30 => sin_inv_data <= to_signed(2,32);
--			when 31 => sin_inv_data <= to_signed(2,32);
--			when 32 => sin_inv_data <= to_signed(2,32);
--			when 33 => sin_inv_data <= to_signed(2,32);
--			when 34 => sin_inv_data <= to_signed(2,32);
--			when 35 => sin_inv_data <= to_signed(2,32);
--			when 36 => sin_inv_data <= to_signed(2,32);
--			when 37 => sin_inv_data <= to_signed(2,32);
--			when 38 => sin_inv_data <= to_signed(2,32);
--			when 39 => sin_inv_data <= to_signed(2,32);
--			when 40 => sin_inv_data <= to_signed(2,32);
--			when 41 => sin_inv_data <= to_signed(2,32);
--			when 42 => sin_inv_data <= to_signed(2,32);
--			when 43 => sin_inv_data <= to_signed(2,32);
--			when 44 => sin_inv_data <= to_signed(3,32);
--			when 45 => sin_inv_data <= to_signed(3,32);
--			when 46 => sin_inv_data <= to_signed(3,32);
--			when 47 => sin_inv_data <= to_signed(3,32);
--			when 48 => sin_inv_data <= to_signed(3,32);
--			when 49 => sin_inv_data <= to_signed(3,32);
--			when 50 => sin_inv_data <= to_signed(3,32);
--			when 51 => sin_inv_data <= to_signed(3,32);
--			when 52 => sin_inv_data <= to_signed(3,32);
--			when 53 => sin_inv_data <= to_signed(3,32);
--			when 54 => sin_inv_data <= to_signed(3,32);
--			when 55 => sin_inv_data <= to_signed(3,32);
--			when 56 => sin_inv_data <= to_signed(3,32);
--			when 57 => sin_inv_data <= to_signed(3,32);
--			when 58 => sin_inv_data <= to_signed(3,32);
--			when 59 => sin_inv_data <= to_signed(3,32);
--			when 60 => sin_inv_data <= to_signed(3,32);
--			when 61 => sin_inv_data <= to_signed(3,32);
--			when 62 => sin_inv_data <= to_signed(4,32);
--			when 63 => sin_inv_data <= to_signed(4,32);
--			when 64 => sin_inv_data <= to_signed(4,32);
--			when 65 => sin_inv_data <= to_signed(4,32);
--			when 66 => sin_inv_data <= to_signed(4,32);
--			when 67 => sin_inv_data <= to_signed(4,32);
--			when 68 => sin_inv_data <= to_signed(4,32);
--			when 69 => sin_inv_data <= to_signed(4,32);
--			when 70 => sin_inv_data <= to_signed(4,32);
--			when 71 => sin_inv_data <= to_signed(4,32);
--			when 72 => sin_inv_data <= to_signed(4,32);
--			when 73 => sin_inv_data <= to_signed(4,32);
--			when 74 => sin_inv_data <= to_signed(4,32);
--			when 75 => sin_inv_data <= to_signed(4,32);
--			when 76 => sin_inv_data <= to_signed(4,32);
--			when 77 => sin_inv_data <= to_signed(4,32);
--			when 78 => sin_inv_data <= to_signed(4,32);
--			when 79 => sin_inv_data <= to_signed(5,32);
--			when 80 => sin_inv_data <= to_signed(5,32);
--			when 81 => sin_inv_data <= to_signed(5,32);
--			when 82 => sin_inv_data <= to_signed(5,32);
--			when 83 => sin_inv_data <= to_signed(5,32);
--			when 84 => sin_inv_data <= to_signed(5,32);
--			when 85 => sin_inv_data <= to_signed(5,32);
--			when 86 => sin_inv_data <= to_signed(5,32);
--			when 87 => sin_inv_data <= to_signed(5,32);
--			when 88 => sin_inv_data <= to_signed(5,32);
--			when 89 => sin_inv_data <= to_signed(5,32);
--			when 90 => sin_inv_data <= to_signed(5,32);
--			when 91 => sin_inv_data <= to_signed(5,32);
--			when 92 => sin_inv_data <= to_signed(5,32);
--			when 93 => sin_inv_data <= to_signed(5,32);
--			when 94 => sin_inv_data <= to_signed(5,32);
--			when 95 => sin_inv_data <= to_signed(5,32);
--			when 96 => sin_inv_data <= to_signed(6,32);
--			when 97 => sin_inv_data <= to_signed(6,32);
--			when 98 => sin_inv_data <= to_signed(6,32);
--			when 99 => sin_inv_data <= to_signed(6,32);
--			when 100 => sin_inv_data <= to_signed(6,32);
--			when 101 => sin_inv_data <= to_signed(6,32);
--			when 102 => sin_inv_data <= to_signed(6,32);
--			when 103 => sin_inv_data <= to_signed(6,32);
--			when 104 => sin_inv_data <= to_signed(6,32);
--			when 105 => sin_inv_data <= to_signed(6,32);
--			when 106 => sin_inv_data <= to_signed(6,32);
--			when 107 => sin_inv_data <= to_signed(6,32);
--			when 108 => sin_inv_data <= to_signed(6,32);
--			when 109 => sin_inv_data <= to_signed(6,32);
--			when 110 => sin_inv_data <= to_signed(6,32);
--			when 111 => sin_inv_data <= to_signed(6,32);
--			when 112 => sin_inv_data <= to_signed(6,32);
--			when 113 => sin_inv_data <= to_signed(6,32);
--			when 114 => sin_inv_data <= to_signed(7,32);
--			when 115 => sin_inv_data <= to_signed(7,32);
--			when 116 => sin_inv_data <= to_signed(7,32);
--			when 117 => sin_inv_data <= to_signed(7,32);
--			when 118 => sin_inv_data <= to_signed(7,32);
--			when 119 => sin_inv_data <= to_signed(7,32);
--			when 120 => sin_inv_data <= to_signed(7,32);
--			when 121 => sin_inv_data <= to_signed(7,32);
--			when 122 => sin_inv_data <= to_signed(7,32);
--			when 123 => sin_inv_data <= to_signed(7,32);
--			when 124 => sin_inv_data <= to_signed(7,32);
--			when 125 => sin_inv_data <= to_signed(7,32);
--			when 126 => sin_inv_data <= to_signed(7,32);
--			when 127 => sin_inv_data <= to_signed(7,32);
--			when 128 => sin_inv_data <= to_signed(7,32);
--			when 129 => sin_inv_data <= to_signed(7,32);
--			when 130 => sin_inv_data <= to_signed(7,32);
--			when 131 => sin_inv_data <= to_signed(8,32);
--			when 132 => sin_inv_data <= to_signed(8,32);
--			when 133 => sin_inv_data <= to_signed(8,32);
--			when 134 => sin_inv_data <= to_signed(8,32);
--			when 135 => sin_inv_data <= to_signed(8,32);
--			when 136 => sin_inv_data <= to_signed(8,32);
--			when 137 => sin_inv_data <= to_signed(8,32);
--			when 138 => sin_inv_data <= to_signed(8,32);
--			when 139 => sin_inv_data <= to_signed(8,32);
--			when 140 => sin_inv_data <= to_signed(8,32);
--			when 141 => sin_inv_data <= to_signed(8,32);
--			when 142 => sin_inv_data <= to_signed(8,32);
--			when 143 => sin_inv_data <= to_signed(8,32);
--			when 144 => sin_inv_data <= to_signed(8,32);
--			when 145 => sin_inv_data <= to_signed(8,32);
--			when 146 => sin_inv_data <= to_signed(8,32);
--			when 147 => sin_inv_data <= to_signed(8,32);
--			when 148 => sin_inv_data <= to_signed(9,32);
--			when 149 => sin_inv_data <= to_signed(9,32);
--			when 150 => sin_inv_data <= to_signed(9,32);
--			when 151 => sin_inv_data <= to_signed(9,32);
--			when 152 => sin_inv_data <= to_signed(9,32);
--			when 153 => sin_inv_data <= to_signed(9,32);
--			when 154 => sin_inv_data <= to_signed(9,32);
--			when 155 => sin_inv_data <= to_signed(9,32);
--			when 156 => sin_inv_data <= to_signed(9,32);
--			when 157 => sin_inv_data <= to_signed(9,32);
--			when 158 => sin_inv_data <= to_signed(9,32);
--			when 159 => sin_inv_data <= to_signed(9,32);
--			when 160 => sin_inv_data <= to_signed(9,32);
--			when 161 => sin_inv_data <= to_signed(9,32);
--			when 162 => sin_inv_data <= to_signed(9,32);
--			when 163 => sin_inv_data <= to_signed(9,32);
--			when 164 => sin_inv_data <= to_signed(9,32);
--			when 165 => sin_inv_data <= to_signed(9,32);
--			when 166 => sin_inv_data <= to_signed(10,32);
--			when 167 => sin_inv_data <= to_signed(10,32);
--			when 168 => sin_inv_data <= to_signed(10,32);
--			when 169 => sin_inv_data <= to_signed(10,32);
--			when 170 => sin_inv_data <= to_signed(10,32);
--			when 171 => sin_inv_data <= to_signed(10,32);
--			when 172 => sin_inv_data <= to_signed(10,32);
--			when 173 => sin_inv_data <= to_signed(10,32);
--			when 174 => sin_inv_data <= to_signed(10,32);
--			when 175 => sin_inv_data <= to_signed(10,32);
--			when 176 => sin_inv_data <= to_signed(10,32);
--			when 177 => sin_inv_data <= to_signed(10,32);
--			when 178 => sin_inv_data <= to_signed(10,32);
--			when 179 => sin_inv_data <= to_signed(10,32);
--			when 180 => sin_inv_data <= to_signed(10,32);
--			when 181 => sin_inv_data <= to_signed(10,32);
--			when 182 => sin_inv_data <= to_signed(10,32);
--			when 183 => sin_inv_data <= to_signed(11,32);
--			when 184 => sin_inv_data <= to_signed(11,32);
--			when 185 => sin_inv_data <= to_signed(11,32);
--			when 186 => sin_inv_data <= to_signed(11,32);
--			when 187 => sin_inv_data <= to_signed(11,32);
--			when 188 => sin_inv_data <= to_signed(11,32);
--			when 189 => sin_inv_data <= to_signed(11,32);
--			when 190 => sin_inv_data <= to_signed(11,32);
--			when 191 => sin_inv_data <= to_signed(11,32);
--			when 192 => sin_inv_data <= to_signed(11,32);
--			when 193 => sin_inv_data <= to_signed(11,32);
--			when 194 => sin_inv_data <= to_signed(11,32);
--			when 195 => sin_inv_data <= to_signed(11,32);
--			when 196 => sin_inv_data <= to_signed(11,32);
--			when 197 => sin_inv_data <= to_signed(11,32);
--			when 198 => sin_inv_data <= to_signed(11,32);
--			when 199 => sin_inv_data <= to_signed(11,32);
--			when 200 => sin_inv_data <= to_signed(12,32);
--			when 201 => sin_inv_data <= to_signed(12,32);
--			when 202 => sin_inv_data <= to_signed(12,32);
--			when 203 => sin_inv_data <= to_signed(12,32);
--			when 204 => sin_inv_data <= to_signed(12,32);
--			when 205 => sin_inv_data <= to_signed(12,32);
--			when 206 => sin_inv_data <= to_signed(12,32);
--			when 207 => sin_inv_data <= to_signed(12,32);
--			when 208 => sin_inv_data <= to_signed(12,32);
--			when 209 => sin_inv_data <= to_signed(12,32);
--			when 210 => sin_inv_data <= to_signed(12,32);
--			when 211 => sin_inv_data <= to_signed(12,32);
--			when 212 => sin_inv_data <= to_signed(12,32);
--			when 213 => sin_inv_data <= to_signed(12,32);
--			when 214 => sin_inv_data <= to_signed(12,32);
--			when 215 => sin_inv_data <= to_signed(12,32);
--			when 216 => sin_inv_data <= to_signed(12,32);
--			when 217 => sin_inv_data <= to_signed(13,32);
--			when 218 => sin_inv_data <= to_signed(13,32);
--			when 219 => sin_inv_data <= to_signed(13,32);
--			when 220 => sin_inv_data <= to_signed(13,32);
--			when 221 => sin_inv_data <= to_signed(13,32);
--			when 222 => sin_inv_data <= to_signed(13,32);
--			when 223 => sin_inv_data <= to_signed(13,32);
--			when 224 => sin_inv_data <= to_signed(13,32);
--			when 225 => sin_inv_data <= to_signed(13,32);
--			when 226 => sin_inv_data <= to_signed(13,32);
--			when 227 => sin_inv_data <= to_signed(13,32);
--			when 228 => sin_inv_data <= to_signed(13,32);
--			when 229 => sin_inv_data <= to_signed(13,32);
--			when 230 => sin_inv_data <= to_signed(13,32);
--			when 231 => sin_inv_data <= to_signed(13,32);
--			when 232 => sin_inv_data <= to_signed(13,32);
--			when 233 => sin_inv_data <= to_signed(13,32);
--			when 234 => sin_inv_data <= to_signed(14,32);
--			when 235 => sin_inv_data <= to_signed(14,32);
--			when 236 => sin_inv_data <= to_signed(14,32);
--			when 237 => sin_inv_data <= to_signed(14,32);
--			when 238 => sin_inv_data <= to_signed(14,32);
--			when 239 => sin_inv_data <= to_signed(14,32);
--			when 240 => sin_inv_data <= to_signed(14,32);
--			when 241 => sin_inv_data <= to_signed(14,32);
--			when 242 => sin_inv_data <= to_signed(14,32);
--			when 243 => sin_inv_data <= to_signed(14,32);
--			when 244 => sin_inv_data <= to_signed(14,32);
--			when 245 => sin_inv_data <= to_signed(14,32);
--			when 246 => sin_inv_data <= to_signed(14,32);
--			when 247 => sin_inv_data <= to_signed(14,32);
--			when 248 => sin_inv_data <= to_signed(14,32);
--			when 249 => sin_inv_data <= to_signed(14,32);
--			when 250 => sin_inv_data <= to_signed(14,32);
--			when 251 => sin_inv_data <= to_signed(15,32);
--			when 252 => sin_inv_data <= to_signed(15,32);
--			when 253 => sin_inv_data <= to_signed(15,32);
--			when 254 => sin_inv_data <= to_signed(15,32);
--			when 255 => sin_inv_data <= to_signed(15,32);
--			when 256 => sin_inv_data <= to_signed(15,32);
--			when 257 => sin_inv_data <= to_signed(15,32);
--			when 258 => sin_inv_data <= to_signed(15,32);
--			when 259 => sin_inv_data <= to_signed(15,32);
--			when 260 => sin_inv_data <= to_signed(15,32);
--			when 261 => sin_inv_data <= to_signed(15,32);
--			when 262 => sin_inv_data <= to_signed(15,32);
--			when 263 => sin_inv_data <= to_signed(15,32);
--			when 264 => sin_inv_data <= to_signed(15,32);
--			when 265 => sin_inv_data <= to_signed(15,32);
--			when 266 => sin_inv_data <= to_signed(15,32);
--			when 267 => sin_inv_data <= to_signed(15,32);
--			when 268 => sin_inv_data <= to_signed(16,32);
--			when 269 => sin_inv_data <= to_signed(16,32);
--			when 270 => sin_inv_data <= to_signed(16,32);
--			when 271 => sin_inv_data <= to_signed(16,32);
--			when 272 => sin_inv_data <= to_signed(16,32);
--			when 273 => sin_inv_data <= to_signed(16,32);
--			when 274 => sin_inv_data <= to_signed(16,32);
--			when 275 => sin_inv_data <= to_signed(16,32);
--			when 276 => sin_inv_data <= to_signed(16,32);
--			when 277 => sin_inv_data <= to_signed(16,32);
--			when 278 => sin_inv_data <= to_signed(16,32);
--			when 279 => sin_inv_data <= to_signed(16,32);
--			when 280 => sin_inv_data <= to_signed(16,32);
--			when 281 => sin_inv_data <= to_signed(16,32);
--			when 282 => sin_inv_data <= to_signed(16,32);
--			when 283 => sin_inv_data <= to_signed(16,32);
--			when 284 => sin_inv_data <= to_signed(16,32);
--			when 285 => sin_inv_data <= to_signed(17,32);
--			when 286 => sin_inv_data <= to_signed(17,32);
--			when 287 => sin_inv_data <= to_signed(17,32);
--			when 288 => sin_inv_data <= to_signed(17,32);
--			when 289 => sin_inv_data <= to_signed(17,32);
--			when 290 => sin_inv_data <= to_signed(17,32);
--			when 291 => sin_inv_data <= to_signed(17,32);
--			when 292 => sin_inv_data <= to_signed(17,32);
--			when 293 => sin_inv_data <= to_signed(17,32);
--			when 294 => sin_inv_data <= to_signed(17,32);
--			when 295 => sin_inv_data <= to_signed(17,32);
--			when 296 => sin_inv_data <= to_signed(17,32);
--			when 297 => sin_inv_data <= to_signed(17,32);
--			when 298 => sin_inv_data <= to_signed(17,32);
--			when 299 => sin_inv_data <= to_signed(17,32);
--			when 300 => sin_inv_data <= to_signed(17,32);
--			when 301 => sin_inv_data <= to_signed(18,32);
--			when 302 => sin_inv_data <= to_signed(18,32);
--			when 303 => sin_inv_data <= to_signed(18,32);
--			when 304 => sin_inv_data <= to_signed(18,32);
--			when 305 => sin_inv_data <= to_signed(18,32);
--			when 306 => sin_inv_data <= to_signed(18,32);
--			when 307 => sin_inv_data <= to_signed(18,32);
--			when 308 => sin_inv_data <= to_signed(18,32);
--			when 309 => sin_inv_data <= to_signed(18,32);
--			when 310 => sin_inv_data <= to_signed(18,32);
--			when 311 => sin_inv_data <= to_signed(18,32);
--			when 312 => sin_inv_data <= to_signed(18,32);
--			when 313 => sin_inv_data <= to_signed(18,32);
--			when 314 => sin_inv_data <= to_signed(18,32);
--			when 315 => sin_inv_data <= to_signed(18,32);
--			when 316 => sin_inv_data <= to_signed(18,32);
--			when 317 => sin_inv_data <= to_signed(18,32);
--			when 318 => sin_inv_data <= to_signed(19,32);
--			when 319 => sin_inv_data <= to_signed(19,32);
--			when 320 => sin_inv_data <= to_signed(19,32);
--			when 321 => sin_inv_data <= to_signed(19,32);
--			when 322 => sin_inv_data <= to_signed(19,32);
--			when 323 => sin_inv_data <= to_signed(19,32);
--			when 324 => sin_inv_data <= to_signed(19,32);
--			when 325 => sin_inv_data <= to_signed(19,32);
--			when 326 => sin_inv_data <= to_signed(19,32);
--			when 327 => sin_inv_data <= to_signed(19,32);
--			when 328 => sin_inv_data <= to_signed(19,32);
--			when 329 => sin_inv_data <= to_signed(19,32);
--			when 330 => sin_inv_data <= to_signed(19,32);
--			when 331 => sin_inv_data <= to_signed(19,32);
--			when 332 => sin_inv_data <= to_signed(19,32);
--			when 333 => sin_inv_data <= to_signed(19,32);
--			when 334 => sin_inv_data <= to_signed(20,32);
--			when 335 => sin_inv_data <= to_signed(20,32);
--			when 336 => sin_inv_data <= to_signed(20,32);
--			when 337 => sin_inv_data <= to_signed(20,32);
--			when 338 => sin_inv_data <= to_signed(20,32);
--			when 339 => sin_inv_data <= to_signed(20,32);
--			when 340 => sin_inv_data <= to_signed(20,32);
--			when 341 => sin_inv_data <= to_signed(20,32);
--			when 342 => sin_inv_data <= to_signed(20,32);
--			when 343 => sin_inv_data <= to_signed(20,32);
--			when 344 => sin_inv_data <= to_signed(20,32);
--			when 345 => sin_inv_data <= to_signed(20,32);
--			when 346 => sin_inv_data <= to_signed(20,32);
--			when 347 => sin_inv_data <= to_signed(20,32);
--			when 348 => sin_inv_data <= to_signed(20,32);
--			when 349 => sin_inv_data <= to_signed(20,32);
--			when 350 => sin_inv_data <= to_signed(20,32);
--			when 351 => sin_inv_data <= to_signed(21,32);
--			when 352 => sin_inv_data <= to_signed(21,32);
--			when 353 => sin_inv_data <= to_signed(21,32);
--			when 354 => sin_inv_data <= to_signed(21,32);
--			when 355 => sin_inv_data <= to_signed(21,32);
--			when 356 => sin_inv_data <= to_signed(21,32);
--			when 357 => sin_inv_data <= to_signed(21,32);
--			when 358 => sin_inv_data <= to_signed(21,32);
--			when 359 => sin_inv_data <= to_signed(21,32);
--			when 360 => sin_inv_data <= to_signed(21,32);
--			when 361 => sin_inv_data <= to_signed(21,32);
--			when 362 => sin_inv_data <= to_signed(21,32);
--			when 363 => sin_inv_data <= to_signed(21,32);
--			when 364 => sin_inv_data <= to_signed(21,32);
--			when 365 => sin_inv_data <= to_signed(21,32);
--			when 366 => sin_inv_data <= to_signed(21,32);
--			when 367 => sin_inv_data <= to_signed(22,32);
--			when 368 => sin_inv_data <= to_signed(22,32);
--			when 369 => sin_inv_data <= to_signed(22,32);
--			when 370 => sin_inv_data <= to_signed(22,32);
--			when 371 => sin_inv_data <= to_signed(22,32);
--			when 372 => sin_inv_data <= to_signed(22,32);
--			when 373 => sin_inv_data <= to_signed(22,32);
--			when 374 => sin_inv_data <= to_signed(22,32);
--			when 375 => sin_inv_data <= to_signed(22,32);
--			when 376 => sin_inv_data <= to_signed(22,32);
--			when 377 => sin_inv_data <= to_signed(22,32);
--			when 378 => sin_inv_data <= to_signed(22,32);
--			when 379 => sin_inv_data <= to_signed(22,32);
--			when 380 => sin_inv_data <= to_signed(22,32);
--			when 381 => sin_inv_data <= to_signed(22,32);
--			when 382 => sin_inv_data <= to_signed(22,32);
--			when 383 => sin_inv_data <= to_signed(23,32);
--			when 384 => sin_inv_data <= to_signed(23,32);
--			when 385 => sin_inv_data <= to_signed(23,32);
--			when 386 => sin_inv_data <= to_signed(23,32);
--			when 387 => sin_inv_data <= to_signed(23,32);
--			when 388 => sin_inv_data <= to_signed(23,32);
--			when 389 => sin_inv_data <= to_signed(23,32);
--			when 390 => sin_inv_data <= to_signed(23,32);
--			when 391 => sin_inv_data <= to_signed(23,32);
--			when 392 => sin_inv_data <= to_signed(23,32);
--			when 393 => sin_inv_data <= to_signed(23,32);
--			when 394 => sin_inv_data <= to_signed(23,32);
--			when 395 => sin_inv_data <= to_signed(23,32);
--			when 396 => sin_inv_data <= to_signed(23,32);
--			when 397 => sin_inv_data <= to_signed(23,32);
--			when 398 => sin_inv_data <= to_signed(23,32);
--			when 399 => sin_inv_data <= to_signed(24,32);
--			when 400 => sin_inv_data <= to_signed(24,32);
--			when 401 => sin_inv_data <= to_signed(24,32);
--			when 402 => sin_inv_data <= to_signed(24,32);
--			when 403 => sin_inv_data <= to_signed(24,32);
--			when 404 => sin_inv_data <= to_signed(24,32);
--			when 405 => sin_inv_data <= to_signed(24,32);
--			when 406 => sin_inv_data <= to_signed(24,32);
--			when 407 => sin_inv_data <= to_signed(24,32);
--			when 408 => sin_inv_data <= to_signed(24,32);
--			when 409 => sin_inv_data <= to_signed(24,32);
--			when 410 => sin_inv_data <= to_signed(24,32);
--			when 411 => sin_inv_data <= to_signed(24,32);
--			when 412 => sin_inv_data <= to_signed(24,32);
--			when 413 => sin_inv_data <= to_signed(24,32);
--			when 414 => sin_inv_data <= to_signed(24,32);
--			when 415 => sin_inv_data <= to_signed(25,32);
--			when 416 => sin_inv_data <= to_signed(25,32);
--			when 417 => sin_inv_data <= to_signed(25,32);
--			when 418 => sin_inv_data <= to_signed(25,32);
--			when 419 => sin_inv_data <= to_signed(25,32);
--			when 420 => sin_inv_data <= to_signed(25,32);
--			when 421 => sin_inv_data <= to_signed(25,32);
--			when 422 => sin_inv_data <= to_signed(25,32);
--			when 423 => sin_inv_data <= to_signed(25,32);
--			when 424 => sin_inv_data <= to_signed(25,32);
--			when 425 => sin_inv_data <= to_signed(25,32);
--			when 426 => sin_inv_data <= to_signed(25,32);
--			when 427 => sin_inv_data <= to_signed(25,32);
--			when 428 => sin_inv_data <= to_signed(25,32);
--			when 429 => sin_inv_data <= to_signed(25,32);
--			when 430 => sin_inv_data <= to_signed(25,32);
--			when 431 => sin_inv_data <= to_signed(26,32);
--			when 432 => sin_inv_data <= to_signed(26,32);
--			when 433 => sin_inv_data <= to_signed(26,32);
--			when 434 => sin_inv_data <= to_signed(26,32);
--			when 435 => sin_inv_data <= to_signed(26,32);
--			when 436 => sin_inv_data <= to_signed(26,32);
--			when 437 => sin_inv_data <= to_signed(26,32);
--			when 438 => sin_inv_data <= to_signed(26,32);
--			when 439 => sin_inv_data <= to_signed(26,32);
--			when 440 => sin_inv_data <= to_signed(26,32);
--			when 441 => sin_inv_data <= to_signed(26,32);
--			when 442 => sin_inv_data <= to_signed(26,32);
--			when 443 => sin_inv_data <= to_signed(26,32);
--			when 444 => sin_inv_data <= to_signed(26,32);
--			when 445 => sin_inv_data <= to_signed(26,32);
--			when 446 => sin_inv_data <= to_signed(26,32);
--			when 447 => sin_inv_data <= to_signed(27,32);
--			when 448 => sin_inv_data <= to_signed(27,32);
--			when 449 => sin_inv_data <= to_signed(27,32);
--			when 450 => sin_inv_data <= to_signed(27,32);
--			when 451 => sin_inv_data <= to_signed(27,32);
--			when 452 => sin_inv_data <= to_signed(27,32);
--			when 453 => sin_inv_data <= to_signed(27,32);
--			when 454 => sin_inv_data <= to_signed(27,32);
--			when 455 => sin_inv_data <= to_signed(27,32);
--			when 456 => sin_inv_data <= to_signed(27,32);
--			when 457 => sin_inv_data <= to_signed(27,32);
--			when 458 => sin_inv_data <= to_signed(27,32);
--			when 459 => sin_inv_data <= to_signed(27,32);
--			when 460 => sin_inv_data <= to_signed(27,32);
--			when 461 => sin_inv_data <= to_signed(27,32);
--			when 462 => sin_inv_data <= to_signed(28,32);
--			when 463 => sin_inv_data <= to_signed(28,32);
--			when 464 => sin_inv_data <= to_signed(28,32);
--			when 465 => sin_inv_data <= to_signed(28,32);
--			when 466 => sin_inv_data <= to_signed(28,32);
--			when 467 => sin_inv_data <= to_signed(28,32);
--			when 468 => sin_inv_data <= to_signed(28,32);
--			when 469 => sin_inv_data <= to_signed(28,32);
--			when 470 => sin_inv_data <= to_signed(28,32);
--			when 471 => sin_inv_data <= to_signed(28,32);
--			when 472 => sin_inv_data <= to_signed(28,32);
--			when 473 => sin_inv_data <= to_signed(28,32);
--			when 474 => sin_inv_data <= to_signed(28,32);
--			when 475 => sin_inv_data <= to_signed(28,32);
--			when 476 => sin_inv_data <= to_signed(28,32);
--			when 477 => sin_inv_data <= to_signed(28,32);
--			when 478 => sin_inv_data <= to_signed(29,32);
--			when 479 => sin_inv_data <= to_signed(29,32);
--			when 480 => sin_inv_data <= to_signed(29,32);
--			when 481 => sin_inv_data <= to_signed(29,32);
--			when 482 => sin_inv_data <= to_signed(29,32);
--			when 483 => sin_inv_data <= to_signed(29,32);
--			when 484 => sin_inv_data <= to_signed(29,32);
--			when 485 => sin_inv_data <= to_signed(29,32);
--			when 486 => sin_inv_data <= to_signed(29,32);
--			when 487 => sin_inv_data <= to_signed(29,32);
--			when 488 => sin_inv_data <= to_signed(29,32);
--			when 489 => sin_inv_data <= to_signed(29,32);
--			when 490 => sin_inv_data <= to_signed(29,32);
--			when 491 => sin_inv_data <= to_signed(29,32);
--			when 492 => sin_inv_data <= to_signed(29,32);
--			when 493 => sin_inv_data <= to_signed(30,32);
--			when 494 => sin_inv_data <= to_signed(30,32);
--			when 495 => sin_inv_data <= to_signed(30,32);
--			when 496 => sin_inv_data <= to_signed(30,32);
--			when 497 => sin_inv_data <= to_signed(30,32);
--			when 498 => sin_inv_data <= to_signed(30,32);
--			when 499 => sin_inv_data <= to_signed(30,32);
--			when 500 => sin_inv_data <= to_signed(30,32);
--			when 501 => sin_inv_data <= to_signed(30,32);
--			when 502 => sin_inv_data <= to_signed(30,32);
--			when 503 => sin_inv_data <= to_signed(30,32);
--			when 504 => sin_inv_data <= to_signed(30,32);
--			when 505 => sin_inv_data <= to_signed(30,32);
--			when 506 => sin_inv_data <= to_signed(30,32);
--			when 507 => sin_inv_data <= to_signed(30,32);
--			when 508 => sin_inv_data <= to_signed(31,32);
--			when 509 => sin_inv_data <= to_signed(31,32);
--			when 510 => sin_inv_data <= to_signed(31,32);
--			when 511 => sin_inv_data <= to_signed(31,32);
--			when 512 => sin_inv_data <= to_signed(31,32);
--			when 513 => sin_inv_data <= to_signed(31,32);
--			when 514 => sin_inv_data <= to_signed(31,32);
--			when 515 => sin_inv_data <= to_signed(31,32);
--			when 516 => sin_inv_data <= to_signed(31,32);
--			when 517 => sin_inv_data <= to_signed(31,32);
--			when 518 => sin_inv_data <= to_signed(31,32);
--			when 519 => sin_inv_data <= to_signed(31,32);
--			when 520 => sin_inv_data <= to_signed(31,32);
--			when 521 => sin_inv_data <= to_signed(31,32);
--			when 522 => sin_inv_data <= to_signed(31,32);
--			when 523 => sin_inv_data <= to_signed(32,32);
--			when 524 => sin_inv_data <= to_signed(32,32);
--			when 525 => sin_inv_data <= to_signed(32,32);
--			when 526 => sin_inv_data <= to_signed(32,32);
--			when 527 => sin_inv_data <= to_signed(32,32);
--			when 528 => sin_inv_data <= to_signed(32,32);
--			when 529 => sin_inv_data <= to_signed(32,32);
--			when 530 => sin_inv_data <= to_signed(32,32);
--			when 531 => sin_inv_data <= to_signed(32,32);
--			when 532 => sin_inv_data <= to_signed(32,32);
--			when 533 => sin_inv_data <= to_signed(32,32);
--			when 534 => sin_inv_data <= to_signed(32,32);
--			when 535 => sin_inv_data <= to_signed(32,32);
--			when 536 => sin_inv_data <= to_signed(32,32);
--			when 537 => sin_inv_data <= to_signed(32,32);
--			when 538 => sin_inv_data <= to_signed(33,32);
--			when 539 => sin_inv_data <= to_signed(33,32);
--			when 540 => sin_inv_data <= to_signed(33,32);
--			when 541 => sin_inv_data <= to_signed(33,32);
--			when 542 => sin_inv_data <= to_signed(33,32);
--			when 543 => sin_inv_data <= to_signed(33,32);
--			when 544 => sin_inv_data <= to_signed(33,32);
--			when 545 => sin_inv_data <= to_signed(33,32);
--			when 546 => sin_inv_data <= to_signed(33,32);
--			when 547 => sin_inv_data <= to_signed(33,32);
--			when 548 => sin_inv_data <= to_signed(33,32);
--			when 549 => sin_inv_data <= to_signed(33,32);
--			when 550 => sin_inv_data <= to_signed(33,32);
--			when 551 => sin_inv_data <= to_signed(33,32);
--			when 552 => sin_inv_data <= to_signed(34,32);
--			when 553 => sin_inv_data <= to_signed(34,32);
--			when 554 => sin_inv_data <= to_signed(34,32);
--			when 555 => sin_inv_data <= to_signed(34,32);
--			when 556 => sin_inv_data <= to_signed(34,32);
--			when 557 => sin_inv_data <= to_signed(34,32);
--			when 558 => sin_inv_data <= to_signed(34,32);
--			when 559 => sin_inv_data <= to_signed(34,32);
--			when 560 => sin_inv_data <= to_signed(34,32);
--			when 561 => sin_inv_data <= to_signed(34,32);
--			when 562 => sin_inv_data <= to_signed(34,32);
--			when 563 => sin_inv_data <= to_signed(34,32);
--			when 564 => sin_inv_data <= to_signed(34,32);
--			when 565 => sin_inv_data <= to_signed(34,32);
--			when 566 => sin_inv_data <= to_signed(34,32);
--			when 567 => sin_inv_data <= to_signed(35,32);
--			when 568 => sin_inv_data <= to_signed(35,32);
--			when 569 => sin_inv_data <= to_signed(35,32);
--			when 570 => sin_inv_data <= to_signed(35,32);
--			when 571 => sin_inv_data <= to_signed(35,32);
--			when 572 => sin_inv_data <= to_signed(35,32);
--			when 573 => sin_inv_data <= to_signed(35,32);
--			when 574 => sin_inv_data <= to_signed(35,32);
--			when 575 => sin_inv_data <= to_signed(35,32);
--			when 576 => sin_inv_data <= to_signed(35,32);
--			when 577 => sin_inv_data <= to_signed(35,32);
--			when 578 => sin_inv_data <= to_signed(35,32);
--			when 579 => sin_inv_data <= to_signed(35,32);
--			when 580 => sin_inv_data <= to_signed(35,32);
--			when 581 => sin_inv_data <= to_signed(36,32);
--			when 582 => sin_inv_data <= to_signed(36,32);
--			when 583 => sin_inv_data <= to_signed(36,32);
--			when 584 => sin_inv_data <= to_signed(36,32);
--			when 585 => sin_inv_data <= to_signed(36,32);
--			when 586 => sin_inv_data <= to_signed(36,32);
--			when 587 => sin_inv_data <= to_signed(36,32);
--			when 588 => sin_inv_data <= to_signed(36,32);
--			when 589 => sin_inv_data <= to_signed(36,32);
--			when 590 => sin_inv_data <= to_signed(36,32);
--			when 591 => sin_inv_data <= to_signed(36,32);
--			when 592 => sin_inv_data <= to_signed(36,32);
--			when 593 => sin_inv_data <= to_signed(36,32);
--			when 594 => sin_inv_data <= to_signed(36,32);
--			when 595 => sin_inv_data <= to_signed(37,32);
--			when 596 => sin_inv_data <= to_signed(37,32);
--			when 597 => sin_inv_data <= to_signed(37,32);
--			when 598 => sin_inv_data <= to_signed(37,32);
--			when 599 => sin_inv_data <= to_signed(37,32);
--			when 600 => sin_inv_data <= to_signed(37,32);
--			when 601 => sin_inv_data <= to_signed(37,32);
--			when 602 => sin_inv_data <= to_signed(37,32);
--			when 603 => sin_inv_data <= to_signed(37,32);
--			when 604 => sin_inv_data <= to_signed(37,32);
--			when 605 => sin_inv_data <= to_signed(37,32);
--			when 606 => sin_inv_data <= to_signed(37,32);
--			when 607 => sin_inv_data <= to_signed(37,32);
--			when 608 => sin_inv_data <= to_signed(37,32);
--			when 609 => sin_inv_data <= to_signed(38,32);
--			when 610 => sin_inv_data <= to_signed(38,32);
--			when 611 => sin_inv_data <= to_signed(38,32);
--			when 612 => sin_inv_data <= to_signed(38,32);
--			when 613 => sin_inv_data <= to_signed(38,32);
--			when 614 => sin_inv_data <= to_signed(38,32);
--			when 615 => sin_inv_data <= to_signed(38,32);
--			when 616 => sin_inv_data <= to_signed(38,32);
--			when 617 => sin_inv_data <= to_signed(38,32);
--			when 618 => sin_inv_data <= to_signed(38,32);
--			when 619 => sin_inv_data <= to_signed(38,32);
--			when 620 => sin_inv_data <= to_signed(38,32);
--			when 621 => sin_inv_data <= to_signed(38,32);
--			when 622 => sin_inv_data <= to_signed(38,32);
--			when 623 => sin_inv_data <= to_signed(39,32);
--			when 624 => sin_inv_data <= to_signed(39,32);
--			when 625 => sin_inv_data <= to_signed(39,32);
--			when 626 => sin_inv_data <= to_signed(39,32);
--			when 627 => sin_inv_data <= to_signed(39,32);
--			when 628 => sin_inv_data <= to_signed(39,32);
--			when 629 => sin_inv_data <= to_signed(39,32);
--			when 630 => sin_inv_data <= to_signed(39,32);
--			when 631 => sin_inv_data <= to_signed(39,32);
--			when 632 => sin_inv_data <= to_signed(39,32);
--			when 633 => sin_inv_data <= to_signed(39,32);
--			when 634 => sin_inv_data <= to_signed(39,32);
--			when 635 => sin_inv_data <= to_signed(39,32);
--			when 636 => sin_inv_data <= to_signed(39,32);
--			when 637 => sin_inv_data <= to_signed(40,32);
--			when 638 => sin_inv_data <= to_signed(40,32);
--			when 639 => sin_inv_data <= to_signed(40,32);
--			when 640 => sin_inv_data <= to_signed(40,32);
--			when 641 => sin_inv_data <= to_signed(40,32);
--			when 642 => sin_inv_data <= to_signed(40,32);
--			when 643 => sin_inv_data <= to_signed(40,32);
--			when 644 => sin_inv_data <= to_signed(40,32);
--			when 645 => sin_inv_data <= to_signed(40,32);
--			when 646 => sin_inv_data <= to_signed(40,32);
--			when 647 => sin_inv_data <= to_signed(40,32);
--			when 648 => sin_inv_data <= to_signed(40,32);
--			when 649 => sin_inv_data <= to_signed(40,32);
--			when 650 => sin_inv_data <= to_signed(41,32);
--			when 651 => sin_inv_data <= to_signed(41,32);
--			when 652 => sin_inv_data <= to_signed(41,32);
--			when 653 => sin_inv_data <= to_signed(41,32);
--			when 654 => sin_inv_data <= to_signed(41,32);
--			when 655 => sin_inv_data <= to_signed(41,32);
--			when 656 => sin_inv_data <= to_signed(41,32);
--			when 657 => sin_inv_data <= to_signed(41,32);
--			when 658 => sin_inv_data <= to_signed(41,32);
--			when 659 => sin_inv_data <= to_signed(41,32);
--			when 660 => sin_inv_data <= to_signed(41,32);
--			when 661 => sin_inv_data <= to_signed(41,32);
--			when 662 => sin_inv_data <= to_signed(41,32);
--			when 663 => sin_inv_data <= to_signed(42,32);
--			when 664 => sin_inv_data <= to_signed(42,32);
--			when 665 => sin_inv_data <= to_signed(42,32);
--			when 666 => sin_inv_data <= to_signed(42,32);
--			when 667 => sin_inv_data <= to_signed(42,32);
--			when 668 => sin_inv_data <= to_signed(42,32);
--			when 669 => sin_inv_data <= to_signed(42,32);
--			when 670 => sin_inv_data <= to_signed(42,32);
--			when 671 => sin_inv_data <= to_signed(42,32);
--			when 672 => sin_inv_data <= to_signed(42,32);
--			when 673 => sin_inv_data <= to_signed(42,32);
--			when 674 => sin_inv_data <= to_signed(42,32);
--			when 675 => sin_inv_data <= to_signed(42,32);
--			when 676 => sin_inv_data <= to_signed(43,32);
--			when 677 => sin_inv_data <= to_signed(43,32);
--			when 678 => sin_inv_data <= to_signed(43,32);
--			when 679 => sin_inv_data <= to_signed(43,32);
--			when 680 => sin_inv_data <= to_signed(43,32);
--			when 681 => sin_inv_data <= to_signed(43,32);
--			when 682 => sin_inv_data <= to_signed(43,32);
--			when 683 => sin_inv_data <= to_signed(43,32);
--			when 684 => sin_inv_data <= to_signed(43,32);
--			when 685 => sin_inv_data <= to_signed(43,32);
--			when 686 => sin_inv_data <= to_signed(43,32);
--			when 687 => sin_inv_data <= to_signed(43,32);
--			when 688 => sin_inv_data <= to_signed(43,32);
--			when 689 => sin_inv_data <= to_signed(44,32);
--			when 690 => sin_inv_data <= to_signed(44,32);
--			when 691 => sin_inv_data <= to_signed(44,32);
--			when 692 => sin_inv_data <= to_signed(44,32);
--			when 693 => sin_inv_data <= to_signed(44,32);
--			when 694 => sin_inv_data <= to_signed(44,32);
--			when 695 => sin_inv_data <= to_signed(44,32);
--			when 696 => sin_inv_data <= to_signed(44,32);
--			when 697 => sin_inv_data <= to_signed(44,32);
--			when 698 => sin_inv_data <= to_signed(44,32);
--			when 699 => sin_inv_data <= to_signed(44,32);
--			when 700 => sin_inv_data <= to_signed(44,32);
--			when 701 => sin_inv_data <= to_signed(45,32);
--			when 702 => sin_inv_data <= to_signed(45,32);
--			when 703 => sin_inv_data <= to_signed(45,32);
--			when 704 => sin_inv_data <= to_signed(45,32);
--			when 705 => sin_inv_data <= to_signed(45,32);
--			when 706 => sin_inv_data <= to_signed(45,32);
--			when 707 => sin_inv_data <= to_signed(45,32);
--			when 708 => sin_inv_data <= to_signed(45,32);
--			when 709 => sin_inv_data <= to_signed(45,32);
--			when 710 => sin_inv_data <= to_signed(45,32);
--			when 711 => sin_inv_data <= to_signed(45,32);
--			when 712 => sin_inv_data <= to_signed(45,32);
--			when 713 => sin_inv_data <= to_signed(45,32);
--			when 714 => sin_inv_data <= to_signed(46,32);
--			when 715 => sin_inv_data <= to_signed(46,32);
--			when 716 => sin_inv_data <= to_signed(46,32);
--			when 717 => sin_inv_data <= to_signed(46,32);
--			when 718 => sin_inv_data <= to_signed(46,32);
--			when 719 => sin_inv_data <= to_signed(46,32);
--			when 720 => sin_inv_data <= to_signed(46,32);
--			when 721 => sin_inv_data <= to_signed(46,32);
--			when 722 => sin_inv_data <= to_signed(46,32);
--			when 723 => sin_inv_data <= to_signed(46,32);
--			when 724 => sin_inv_data <= to_signed(46,32);
--			when 725 => sin_inv_data <= to_signed(46,32);
--			when 726 => sin_inv_data <= to_signed(47,32);
--			when 727 => sin_inv_data <= to_signed(47,32);
--			when 728 => sin_inv_data <= to_signed(47,32);
--			when 729 => sin_inv_data <= to_signed(47,32);
--			when 730 => sin_inv_data <= to_signed(47,32);
--			when 731 => sin_inv_data <= to_signed(47,32);
--			when 732 => sin_inv_data <= to_signed(47,32);
--			when 733 => sin_inv_data <= to_signed(47,32);
--			when 734 => sin_inv_data <= to_signed(47,32);
--			when 735 => sin_inv_data <= to_signed(47,32);
--			when 736 => sin_inv_data <= to_signed(47,32);
--			when 737 => sin_inv_data <= to_signed(47,32);
--			when 738 => sin_inv_data <= to_signed(48,32);
--			when 739 => sin_inv_data <= to_signed(48,32);
--			when 740 => sin_inv_data <= to_signed(48,32);
--			when 741 => sin_inv_data <= to_signed(48,32);
--			when 742 => sin_inv_data <= to_signed(48,32);
--			when 743 => sin_inv_data <= to_signed(48,32);
--			when 744 => sin_inv_data <= to_signed(48,32);
--			when 745 => sin_inv_data <= to_signed(48,32);
--			when 746 => sin_inv_data <= to_signed(48,32);
--			when 747 => sin_inv_data <= to_signed(48,32);
--			when 748 => sin_inv_data <= to_signed(48,32);
--			when 749 => sin_inv_data <= to_signed(49,32);
--			when 750 => sin_inv_data <= to_signed(49,32);
--			when 751 => sin_inv_data <= to_signed(49,32);
--			when 752 => sin_inv_data <= to_signed(49,32);
--			when 753 => sin_inv_data <= to_signed(49,32);
--			when 754 => sin_inv_data <= to_signed(49,32);
--			when 755 => sin_inv_data <= to_signed(49,32);
--			when 756 => sin_inv_data <= to_signed(49,32);
--			when 757 => sin_inv_data <= to_signed(49,32);
--			when 758 => sin_inv_data <= to_signed(49,32);
--			when 759 => sin_inv_data <= to_signed(49,32);
--			when 760 => sin_inv_data <= to_signed(49,32);
--			when 761 => sin_inv_data <= to_signed(50,32);
--			when 762 => sin_inv_data <= to_signed(50,32);
--			when 763 => sin_inv_data <= to_signed(50,32);
--			when 764 => sin_inv_data <= to_signed(50,32);
--			when 765 => sin_inv_data <= to_signed(50,32);
--			when 766 => sin_inv_data <= to_signed(50,32);
--			when 767 => sin_inv_data <= to_signed(50,32);
--			when 768 => sin_inv_data <= to_signed(50,32);
--			when 769 => sin_inv_data <= to_signed(50,32);
--			when 770 => sin_inv_data <= to_signed(50,32);
--			when 771 => sin_inv_data <= to_signed(50,32);
--			when 772 => sin_inv_data <= to_signed(51,32);
--			when 773 => sin_inv_data <= to_signed(51,32);
--			when 774 => sin_inv_data <= to_signed(51,32);
--			when 775 => sin_inv_data <= to_signed(51,32);
--			when 776 => sin_inv_data <= to_signed(51,32);
--			when 777 => sin_inv_data <= to_signed(51,32);
--			when 778 => sin_inv_data <= to_signed(51,32);
--			when 779 => sin_inv_data <= to_signed(51,32);
--			when 780 => sin_inv_data <= to_signed(51,32);
--			when 781 => sin_inv_data <= to_signed(51,32);
--			when 782 => sin_inv_data <= to_signed(51,32);
--			when 783 => sin_inv_data <= to_signed(52,32);
--			when 784 => sin_inv_data <= to_signed(52,32);
--			when 785 => sin_inv_data <= to_signed(52,32);
--			when 786 => sin_inv_data <= to_signed(52,32);
--			when 787 => sin_inv_data <= to_signed(52,32);
--			when 788 => sin_inv_data <= to_signed(52,32);
--			when 789 => sin_inv_data <= to_signed(52,32);
--			when 790 => sin_inv_data <= to_signed(52,32);
--			when 791 => sin_inv_data <= to_signed(52,32);
--			when 792 => sin_inv_data <= to_signed(52,32);
--			when 793 => sin_inv_data <= to_signed(52,32);
--			when 794 => sin_inv_data <= to_signed(53,32);
--			when 795 => sin_inv_data <= to_signed(53,32);
--			when 796 => sin_inv_data <= to_signed(53,32);
--			when 797 => sin_inv_data <= to_signed(53,32);
--			when 798 => sin_inv_data <= to_signed(53,32);
--			when 799 => sin_inv_data <= to_signed(53,32);
--			when 800 => sin_inv_data <= to_signed(53,32);
--			when 801 => sin_inv_data <= to_signed(53,32);
--			when 802 => sin_inv_data <= to_signed(53,32);
--			when 803 => sin_inv_data <= to_signed(53,32);
--			when 804 => sin_inv_data <= to_signed(54,32);
--			when 805 => sin_inv_data <= to_signed(54,32);
--			when 806 => sin_inv_data <= to_signed(54,32);
--			when 807 => sin_inv_data <= to_signed(54,32);
--			when 808 => sin_inv_data <= to_signed(54,32);
--			when 809 => sin_inv_data <= to_signed(54,32);
--			when 810 => sin_inv_data <= to_signed(54,32);
--			when 811 => sin_inv_data <= to_signed(54,32);
--			when 812 => sin_inv_data <= to_signed(54,32);
--			when 813 => sin_inv_data <= to_signed(54,32);
--			when 814 => sin_inv_data <= to_signed(54,32);
--			when 815 => sin_inv_data <= to_signed(55,32);
--			when 816 => sin_inv_data <= to_signed(55,32);
--			when 817 => sin_inv_data <= to_signed(55,32);
--			when 818 => sin_inv_data <= to_signed(55,32);
--			when 819 => sin_inv_data <= to_signed(55,32);
--			when 820 => sin_inv_data <= to_signed(55,32);
--			when 821 => sin_inv_data <= to_signed(55,32);
--			when 822 => sin_inv_data <= to_signed(55,32);
--			when 823 => sin_inv_data <= to_signed(55,32);
--			when 824 => sin_inv_data <= to_signed(55,32);
--			when 825 => sin_inv_data <= to_signed(56,32);
--			when 826 => sin_inv_data <= to_signed(56,32);
--			when 827 => sin_inv_data <= to_signed(56,32);
--			when 828 => sin_inv_data <= to_signed(56,32);
--			when 829 => sin_inv_data <= to_signed(56,32);
--			when 830 => sin_inv_data <= to_signed(56,32);
--			when 831 => sin_inv_data <= to_signed(56,32);
--			when 832 => sin_inv_data <= to_signed(56,32);
--			when 833 => sin_inv_data <= to_signed(56,32);
--			when 834 => sin_inv_data <= to_signed(57,32);
--			when 835 => sin_inv_data <= to_signed(57,32);
--			when 836 => sin_inv_data <= to_signed(57,32);
--			when 837 => sin_inv_data <= to_signed(57,32);
--			when 838 => sin_inv_data <= to_signed(57,32);
--			when 839 => sin_inv_data <= to_signed(57,32);
--			when 840 => sin_inv_data <= to_signed(57,32);
--			when 841 => sin_inv_data <= to_signed(57,32);
--			when 842 => sin_inv_data <= to_signed(57,32);
--			when 843 => sin_inv_data <= to_signed(57,32);
--			when 844 => sin_inv_data <= to_signed(58,32);
--			when 845 => sin_inv_data <= to_signed(58,32);
--			when 846 => sin_inv_data <= to_signed(58,32);
--			when 847 => sin_inv_data <= to_signed(58,32);
--			when 848 => sin_inv_data <= to_signed(58,32);
--			when 849 => sin_inv_data <= to_signed(58,32);
--			when 850 => sin_inv_data <= to_signed(58,32);
--			when 851 => sin_inv_data <= to_signed(58,32);
--			when 852 => sin_inv_data <= to_signed(58,32);
--			when 853 => sin_inv_data <= to_signed(59,32);
--			when 854 => sin_inv_data <= to_signed(59,32);
--			when 855 => sin_inv_data <= to_signed(59,32);
--			when 856 => sin_inv_data <= to_signed(59,32);
--			when 857 => sin_inv_data <= to_signed(59,32);
--			when 858 => sin_inv_data <= to_signed(59,32);
--			when 859 => sin_inv_data <= to_signed(59,32);
--			when 860 => sin_inv_data <= to_signed(59,32);
--			when 861 => sin_inv_data <= to_signed(59,32);
--			when 862 => sin_inv_data <= to_signed(60,32);
--			when 863 => sin_inv_data <= to_signed(60,32);
--			when 864 => sin_inv_data <= to_signed(60,32);
--			when 865 => sin_inv_data <= to_signed(60,32);
--			when 866 => sin_inv_data <= to_signed(60,32);
--			when 867 => sin_inv_data <= to_signed(60,32);
--			when 868 => sin_inv_data <= to_signed(60,32);
--			when 869 => sin_inv_data <= to_signed(60,32);
--			when 870 => sin_inv_data <= to_signed(60,32);
--			when 871 => sin_inv_data <= to_signed(61,32);
--			when 872 => sin_inv_data <= to_signed(61,32);
--			when 873 => sin_inv_data <= to_signed(61,32);
--			when 874 => sin_inv_data <= to_signed(61,32);
--			when 875 => sin_inv_data <= to_signed(61,32);
--			when 876 => sin_inv_data <= to_signed(61,32);
--			when 877 => sin_inv_data <= to_signed(61,32);
--			when 878 => sin_inv_data <= to_signed(61,32);
--			when 879 => sin_inv_data <= to_signed(62,32);
--			when 880 => sin_inv_data <= to_signed(62,32);
--			when 881 => sin_inv_data <= to_signed(62,32);
--			when 882 => sin_inv_data <= to_signed(62,32);
--			when 883 => sin_inv_data <= to_signed(62,32);
--			when 884 => sin_inv_data <= to_signed(62,32);
--			when 885 => sin_inv_data <= to_signed(62,32);
--			when 886 => sin_inv_data <= to_signed(62,32);
--			when 887 => sin_inv_data <= to_signed(62,32);
--			when 888 => sin_inv_data <= to_signed(63,32);
--			when 889 => sin_inv_data <= to_signed(63,32);
--			when 890 => sin_inv_data <= to_signed(63,32);
--			when 891 => sin_inv_data <= to_signed(63,32);
--			when 892 => sin_inv_data <= to_signed(63,32);
--			when 893 => sin_inv_data <= to_signed(63,32);
--			when 894 => sin_inv_data <= to_signed(63,32);
--			when 895 => sin_inv_data <= to_signed(64,32);
--			when 896 => sin_inv_data <= to_signed(64,32);
--			when 897 => sin_inv_data <= to_signed(64,32);
--			when 898 => sin_inv_data <= to_signed(64,32);
--			when 899 => sin_inv_data <= to_signed(64,32);
--			when 900 => sin_inv_data <= to_signed(64,32);
--			when 901 => sin_inv_data <= to_signed(64,32);
--			when 902 => sin_inv_data <= to_signed(64,32);
--			when 903 => sin_inv_data <= to_signed(65,32);
--			when 904 => sin_inv_data <= to_signed(65,32);
--			when 905 => sin_inv_data <= to_signed(65,32);
--			when 906 => sin_inv_data <= to_signed(65,32);
--			when 907 => sin_inv_data <= to_signed(65,32);
--			when 908 => sin_inv_data <= to_signed(65,32);
--			when 909 => sin_inv_data <= to_signed(65,32);
--			when 910 => sin_inv_data <= to_signed(66,32);
--			when 911 => sin_inv_data <= to_signed(66,32);
--			when 912 => sin_inv_data <= to_signed(66,32);
--			when 913 => sin_inv_data <= to_signed(66,32);
--			when 914 => sin_inv_data <= to_signed(66,32);
--			when 915 => sin_inv_data <= to_signed(66,32);
--			when 916 => sin_inv_data <= to_signed(66,32);
--			when 917 => sin_inv_data <= to_signed(66,32);
--			when 918 => sin_inv_data <= to_signed(67,32);
--			when 919 => sin_inv_data <= to_signed(67,32);
--			when 920 => sin_inv_data <= to_signed(67,32);
--			when 921 => sin_inv_data <= to_signed(67,32);
--			when 922 => sin_inv_data <= to_signed(67,32);
--			when 923 => sin_inv_data <= to_signed(67,32);
--			when 924 => sin_inv_data <= to_signed(68,32);
--			when 925 => sin_inv_data <= to_signed(68,32);
--			when 926 => sin_inv_data <= to_signed(68,32);
--			when 927 => sin_inv_data <= to_signed(68,32);
--			when 928 => sin_inv_data <= to_signed(68,32);
--			when 929 => sin_inv_data <= to_signed(68,32);
--			when 930 => sin_inv_data <= to_signed(68,32);
--			when 931 => sin_inv_data <= to_signed(69,32);
--			when 932 => sin_inv_data <= to_signed(69,32);
--			when 933 => sin_inv_data <= to_signed(69,32);
--			when 934 => sin_inv_data <= to_signed(69,32);
--			when 935 => sin_inv_data <= to_signed(69,32);
--			when 936 => sin_inv_data <= to_signed(69,32);
--			when 937 => sin_inv_data <= to_signed(70,32);
--			when 938 => sin_inv_data <= to_signed(70,32);
--			when 939 => sin_inv_data <= to_signed(70,32);
--			when 940 => sin_inv_data <= to_signed(70,32);
--			when 941 => sin_inv_data <= to_signed(70,32);
--			when 942 => sin_inv_data <= to_signed(70,32);
--			when 943 => sin_inv_data <= to_signed(71,32);
--			when 944 => sin_inv_data <= to_signed(71,32);
--			when 945 => sin_inv_data <= to_signed(71,32);
--			when 946 => sin_inv_data <= to_signed(71,32);
--			when 947 => sin_inv_data <= to_signed(71,32);
--			when 948 => sin_inv_data <= to_signed(71,32);
--			when 949 => sin_inv_data <= to_signed(72,32);
--			when 950 => sin_inv_data <= to_signed(72,32);
--			when 951 => sin_inv_data <= to_signed(72,32);
--			when 952 => sin_inv_data <= to_signed(72,32);
--			when 953 => sin_inv_data <= to_signed(72,32);
--			when 954 => sin_inv_data <= to_signed(73,32);
--			when 955 => sin_inv_data <= to_signed(73,32);
--			when 956 => sin_inv_data <= to_signed(73,32);
--			when 957 => sin_inv_data <= to_signed(73,32);
--			when 958 => sin_inv_data <= to_signed(73,32);
--			when 959 => sin_inv_data <= to_signed(74,32);
--			when 960 => sin_inv_data <= to_signed(74,32);
--			when 961 => sin_inv_data <= to_signed(74,32);
--			when 962 => sin_inv_data <= to_signed(74,32);
--			when 963 => sin_inv_data <= to_signed(74,32);
--			when 964 => sin_inv_data <= to_signed(75,32);
--			when 965 => sin_inv_data <= to_signed(75,32);
--			when 966 => sin_inv_data <= to_signed(75,32);
--			when 967 => sin_inv_data <= to_signed(75,32);
--			when 968 => sin_inv_data <= to_signed(75,32);
--			when 969 => sin_inv_data <= to_signed(76,32);
--			when 970 => sin_inv_data <= to_signed(76,32);
--			when 971 => sin_inv_data <= to_signed(76,32);
--			when 972 => sin_inv_data <= to_signed(76,32);
--			when 973 => sin_inv_data <= to_signed(77,32);
--			when 974 => sin_inv_data <= to_signed(77,32);
--			when 975 => sin_inv_data <= to_signed(77,32);
--			when 976 => sin_inv_data <= to_signed(77,32);
--			when 977 => sin_inv_data <= to_signed(78,32);
--			when 978 => sin_inv_data <= to_signed(78,32);
--			when 979 => sin_inv_data <= to_signed(78,32);
--			when 980 => sin_inv_data <= to_signed(79,32);
--			when 981 => sin_inv_data <= to_signed(79,32);
--			when 982 => sin_inv_data <= to_signed(79,32);
--			when 983 => sin_inv_data <= to_signed(79,32);
--			when 984 => sin_inv_data <= to_signed(80,32);
--			when 985 => sin_inv_data <= to_signed(80,32);
--			when 986 => sin_inv_data <= to_signed(80,32);
--			when 987 => sin_inv_data <= to_signed(81,32);
--			when 988 => sin_inv_data <= to_signed(81,32);
--			when 989 => sin_inv_data <= to_signed(81,32);
--			when 990 => sin_inv_data <= to_signed(82,32);
--			when 991 => sin_inv_data <= to_signed(82,32);
--			when 992 => sin_inv_data <= to_signed(83,32);
--			when 993 => sin_inv_data <= to_signed(83,32);
--			when 994 => sin_inv_data <= to_signed(84,32);
--			when 995 => sin_inv_data <= to_signed(84,32);
--			when 996 => sin_inv_data <= to_signed(85,32);
--			when 997 => sin_inv_data <= to_signed(86,32);
--			when 998 => sin_inv_data <= to_signed(86,32);
--			when 999 => sin_inv_data <= to_signed(87,32);
--			when 1000 => sin_inv_data <= to_signed(90,32);
--
--      when others       => null;
--      end case;
--
--      
	      case theta_int_inv is
			when -1000 => sin_inv_data <=   -90;
			when -999 => sin_inv_data <=  -87;
			when -998 => sin_inv_data <=  -86;
			when -997 => sin_inv_data <=  -86;
			when -996 => sin_inv_data <=  -85;
			when -995 => sin_inv_data <=  -84;
			when -994 => sin_inv_data <=  -84;
			when -993 => sin_inv_data <=  -83;
			when -992 => sin_inv_data <=  -83;
			when -991 => sin_inv_data <=  -82;
			when -990 => sin_inv_data <=  -82;
			when -989 => sin_inv_data <=  -81;
			when -988 => sin_inv_data <=  -81;
			when -987 => sin_inv_data <=  -81;
			when -986 => sin_inv_data <=  -80;
			when -985 => sin_inv_data <=  -80;
			when -984 => sin_inv_data <=  -80;
			when -983 => sin_inv_data <=  -79;
			when -982 => sin_inv_data <=  -79;
			when -981 => sin_inv_data <=  -79;
			when -980 => sin_inv_data <=  -79;
			when -979 => sin_inv_data <=  -78;
			when -978 => sin_inv_data <=  -78;
			when -977 => sin_inv_data <=  -78;
			when -976 => sin_inv_data <=  -77;
			when -975 => sin_inv_data <=  -77;
			when -974 => sin_inv_data <=  -77;
			when -973 => sin_inv_data <=  -77;
			when -972 => sin_inv_data <=  -76;
			when -971 => sin_inv_data <=  -76;
			when -970 => sin_inv_data <=  -76;
			when -969 => sin_inv_data <=  -76;
			when -968 => sin_inv_data <=  -75;
			when -967 => sin_inv_data <=  -75;
			when -966 => sin_inv_data <=  -75;
			when -965 => sin_inv_data <=  -75;
			when -964 => sin_inv_data <=  -75;
			when -963 => sin_inv_data <=  -74;
			when -962 => sin_inv_data <=  -74;
			when -961 => sin_inv_data <=  -74;
			when -960 => sin_inv_data <=  -74;
			when -959 => sin_inv_data <=  -74;
			when -958 => sin_inv_data <=  -73;
			when -957 => sin_inv_data <=  -73;
			when -956 => sin_inv_data <=  -73;
			when -955 => sin_inv_data <=  -73;
			when -954 => sin_inv_data <=  -73;
			when -953 => sin_inv_data <=  -72;
			when -952 => sin_inv_data <=  -72;
			when -951 => sin_inv_data <=  -72;
			when -950 => sin_inv_data <=  -72;
			when -949 => sin_inv_data <=  -72;
			when -948 => sin_inv_data <=  -71;
			when -947 => sin_inv_data <=  -71;
			when -946 => sin_inv_data <=  -71;
			when -945 => sin_inv_data <=  -71;
			when -944 => sin_inv_data <=  -71;
			when -943 => sin_inv_data <=  -71;
			when -942 => sin_inv_data <=  -70;
			when -941 => sin_inv_data <=  -70;
			when -940 => sin_inv_data <=  -70;
			when -939 => sin_inv_data <=  -70;
			when -938 => sin_inv_data <=  -70;
			when -937 => sin_inv_data <=  -70;
			when -936 => sin_inv_data <=  -69;
			when -935 => sin_inv_data <=  -69;
			when -934 => sin_inv_data <=  -69;
			when -933 => sin_inv_data <=  -69;
			when -932 => sin_inv_data <=  -69;
			when -931 => sin_inv_data <=  -69;
			when -930 => sin_inv_data <=  -68;
			when -929 => sin_inv_data <=  -68;
			when -928 => sin_inv_data <=  -68;
			when -927 => sin_inv_data <=  -68;
			when -926 => sin_inv_data <=  -68;
			when -925 => sin_inv_data <=  -68;
			when -924 => sin_inv_data <=  -68;
			when -923 => sin_inv_data <=  -67;
			when -922 => sin_inv_data <=  -67;
			when -921 => sin_inv_data <=  -67;
			when -920 => sin_inv_data <=  -67;
			when -919 => sin_inv_data <=  -67;
			when -918 => sin_inv_data <=  -67;
			when -917 => sin_inv_data <=  -66;
			when -916 => sin_inv_data <=  -66;
			when -915 => sin_inv_data <=  -66;
			when -914 => sin_inv_data <=  -66;
			when -913 => sin_inv_data <=  -66;
			when -912 => sin_inv_data <=  -66;
			when -911 => sin_inv_data <=  -66;
			when -910 => sin_inv_data <=  -66;
			when -909 => sin_inv_data <=  -65;
			when -908 => sin_inv_data <=  -65;
			when -907 => sin_inv_data <=  -65;
			when -906 => sin_inv_data <=  -65;
			when -905 => sin_inv_data <=  -65;
			when -904 => sin_inv_data <=  -65;
			when -903 => sin_inv_data <=  -65;
			when -902 => sin_inv_data <=  -64;
			when -901 => sin_inv_data <=  -64;
			when -900 => sin_inv_data <=  -64;
			when -899 => sin_inv_data <=  -64;
			when -898 => sin_inv_data <=  -64;
			when -897 => sin_inv_data <=  -64;
			when -896 => sin_inv_data <=  -64;
			when -895 => sin_inv_data <=  -64;
			when -894 => sin_inv_data <=  -63;
			when -893 => sin_inv_data <=  -63;
			when -892 => sin_inv_data <=  -63;
			when -891 => sin_inv_data <=  -63;
			when -890 => sin_inv_data <=  -63;
			when -889 => sin_inv_data <=  -63;
			when -888 => sin_inv_data <=  -63;
			when -887 => sin_inv_data <=  -62;
			when -886 => sin_inv_data <=  -62;
			when -885 => sin_inv_data <=  -62;
			when -884 => sin_inv_data <=  -62;
			when -883 => sin_inv_data <=  -62;
			when -882 => sin_inv_data <=  -62;
			when -881 => sin_inv_data <=  -62;
			when -880 => sin_inv_data <=  -62;
			when -879 => sin_inv_data <=  -62;
			when -878 => sin_inv_data <=  -61;
			when -877 => sin_inv_data <=  -61;
			when -876 => sin_inv_data <=  -61;
			when -875 => sin_inv_data <=  -61;
			when -874 => sin_inv_data <=  -61;
			when -873 => sin_inv_data <=  -61;
			when -872 => sin_inv_data <=  -61;
			when -871 => sin_inv_data <=  -61;
			when -870 => sin_inv_data <=  -60;
			when -869 => sin_inv_data <=  -60;
			when -868 => sin_inv_data <=  -60;
			when -867 => sin_inv_data <=  -60;
			when -866 => sin_inv_data <=  -60;
			when -865 => sin_inv_data <=  -60;
			when -864 => sin_inv_data <=  -60;
			when -863 => sin_inv_data <=  -60;
			when -862 => sin_inv_data <=  -60;
			when -861 => sin_inv_data <=  -59;
			when -860 => sin_inv_data <=  -59;
			when -859 => sin_inv_data <=  -59;
			when -858 => sin_inv_data <=  -59;
			when -857 => sin_inv_data <=  -59;
			when -856 => sin_inv_data <=  -59;
			when -855 => sin_inv_data <=  -59;
			when -854 => sin_inv_data <=  -59;
			when -853 => sin_inv_data <=  -59;
			when -852 => sin_inv_data <=  -58;
			when -851 => sin_inv_data <=  -58;
			when -850 => sin_inv_data <=  -58;
			when -849 => sin_inv_data <=  -58;
			when -848 => sin_inv_data <=  -58;
			when -847 => sin_inv_data <=  -58;
			when -846 => sin_inv_data <=  -58;
			when -845 => sin_inv_data <=  -58;
			when -844 => sin_inv_data <=  -58;
			when -843 => sin_inv_data <=  -57;
			when -842 => sin_inv_data <=  -57;
			when -841 => sin_inv_data <=  -57;
			when -840 => sin_inv_data <=  -57;
			when -839 => sin_inv_data <=  -57;
			when -838 => sin_inv_data <=  -57;
			when -837 => sin_inv_data <=  -57;
			when -836 => sin_inv_data <=  -57;
			when -835 => sin_inv_data <=  -57;
			when -834 => sin_inv_data <=  -57;
			when -833 => sin_inv_data <=  -56;
			when -832 => sin_inv_data <=  -56;
			when -831 => sin_inv_data <=  -56;
			when -830 => sin_inv_data <=  -56;
			when -829 => sin_inv_data <=  -56;
			when -828 => sin_inv_data <=  -56;
			when -827 => sin_inv_data <=  -56;
			when -826 => sin_inv_data <=  -56;
			when -825 => sin_inv_data <=  -56;
			when -824 => sin_inv_data <=  -55;
			when -823 => sin_inv_data <=  -55;
			when -822 => sin_inv_data <=  -55;
			when -821 => sin_inv_data <=  -55;
			when -820 => sin_inv_data <=  -55;
			when -819 => sin_inv_data <=  -55;
			when -818 => sin_inv_data <=  -55;
			when -817 => sin_inv_data <=  -55;
			when -816 => sin_inv_data <=  -55;
			when -815 => sin_inv_data <=  -55;
			when -814 => sin_inv_data <=  -54;
			when -813 => sin_inv_data <=  -54;
			when -812 => sin_inv_data <=  -54;
			when -811 => sin_inv_data <=  -54;
			when -810 => sin_inv_data <=  -54;
			when -809 => sin_inv_data <=  -54;
			when -808 => sin_inv_data <=  -54;
			when -807 => sin_inv_data <=  -54;
			when -806 => sin_inv_data <=  -54;
			when -805 => sin_inv_data <=  -54;
			when -804 => sin_inv_data <=  -54;
			when -803 => sin_inv_data <=  -53;
			when -802 => sin_inv_data <=  -53;
			when -801 => sin_inv_data <=  -53;
			when -800 => sin_inv_data <=  -53;
			when -799 => sin_inv_data <=  -53;
			when -798 => sin_inv_data <=  -53;
			when -797 => sin_inv_data <=  -53;
			when -796 => sin_inv_data <=  -53;
			when -795 => sin_inv_data <=  -53;
			when -794 => sin_inv_data <=  -53;
			when -793 => sin_inv_data <=  -52;
			when -792 => sin_inv_data <=  -52;
			when -791 => sin_inv_data <=  -52;
			when -790 => sin_inv_data <=  -52;
			when -789 => sin_inv_data <=  -52;
			when -788 => sin_inv_data <=  -52;
			when -787 => sin_inv_data <=  -52;
			when -786 => sin_inv_data <=  -52;
			when -785 => sin_inv_data <=  -52;
			when -784 => sin_inv_data <=  -52;
			when -783 => sin_inv_data <=  -52;
			when -782 => sin_inv_data <=  -51;
			when -781 => sin_inv_data <=  -51;
			when -780 => sin_inv_data <=  -51;
			when -779 => sin_inv_data <=  -51;
			when -778 => sin_inv_data <=  -51;
			when -777 => sin_inv_data <=  -51;
			when -776 => sin_inv_data <=  -51;
			when -775 => sin_inv_data <=  -51;
			when -774 => sin_inv_data <=  -51;
			when -773 => sin_inv_data <=  -51;
			when -772 => sin_inv_data <=  -51;
			when -771 => sin_inv_data <=  -50;
			when -770 => sin_inv_data <=  -50;
			when -769 => sin_inv_data <=  -50;
			when -768 => sin_inv_data <=  -50;
			when -767 => sin_inv_data <=  -50;
			when -766 => sin_inv_data <=  -50;
			when -765 => sin_inv_data <=  -50;
			when -764 => sin_inv_data <=  -50;
			when -763 => sin_inv_data <=  -50;
			when -762 => sin_inv_data <=  -50;
			when -761 => sin_inv_data <=  -50;
			when -760 => sin_inv_data <=  -49;
			when -759 => sin_inv_data <=  -49;
			when -758 => sin_inv_data <=  -49;
			when -757 => sin_inv_data <=  -49;
			when -756 => sin_inv_data <=  -49;
			when -755 => sin_inv_data <=  -49;
			when -754 => sin_inv_data <=  -49;
			when -753 => sin_inv_data <=  -49;
			when -752 => sin_inv_data <=  -49;
			when -751 => sin_inv_data <=  -49;
			when -750 => sin_inv_data <=  -49;
			when -749 => sin_inv_data <=  -49;
			when -748 => sin_inv_data <=  -48;
			when -747 => sin_inv_data <=  -48;
			when -746 => sin_inv_data <=  -48;
			when -745 => sin_inv_data <=  -48;
			when -744 => sin_inv_data <=  -48;
			when -743 => sin_inv_data <=  -48;
			when -742 => sin_inv_data <=  -48;
			when -741 => sin_inv_data <=  -48;
			when -740 => sin_inv_data <=  -48;
			when -739 => sin_inv_data <=  -48;
			when -738 => sin_inv_data <=  -48;
			when -737 => sin_inv_data <=  -47;
			when -736 => sin_inv_data <=  -47;
			when -735 => sin_inv_data <=  -47;
			when -734 => sin_inv_data <=  -47;
			when -733 => sin_inv_data <=  -47;
			when -732 => sin_inv_data <=  -47;
			when -731 => sin_inv_data <=  -47;
			when -730 => sin_inv_data <=  -47;
			when -729 => sin_inv_data <=  -47;
			when -728 => sin_inv_data <=  -47;
			when -727 => sin_inv_data <=  -47;
			when -726 => sin_inv_data <=  -47;
			when -725 => sin_inv_data <=  -46;
			when -724 => sin_inv_data <=  -46;
			when -723 => sin_inv_data <=  -46;
			when -722 => sin_inv_data <=  -46;
			when -721 => sin_inv_data <=  -46;
			when -720 => sin_inv_data <=  -46;
			when -719 => sin_inv_data <=  -46;
			when -718 => sin_inv_data <=  -46;
			when -717 => sin_inv_data <=  -46;
			when -716 => sin_inv_data <=  -46;
			when -715 => sin_inv_data <=  -46;
			when -714 => sin_inv_data <=  -46;
			when -713 => sin_inv_data <=  -45;
			when -712 => sin_inv_data <=  -45;
			when -711 => sin_inv_data <=  -45;
			when -710 => sin_inv_data <=  -45;
			when -709 => sin_inv_data <=  -45;
			when -708 => sin_inv_data <=  -45;
			when -707 => sin_inv_data <=  -45;
			when -706 => sin_inv_data <=  -45;
			when -705 => sin_inv_data <=  -45;
			when -704 => sin_inv_data <=  -45;
			when -703 => sin_inv_data <=  -45;
			when -702 => sin_inv_data <=  -45;
			when -701 => sin_inv_data <=  -45;
			when -700 => sin_inv_data <=  -44;
			when -699 => sin_inv_data <=  -44;
			when -698 => sin_inv_data <=  -44;
			when -697 => sin_inv_data <=  -44;
			when -696 => sin_inv_data <=  -44;
			when -695 => sin_inv_data <=  -44;
			when -694 => sin_inv_data <=  -44;
			when -693 => sin_inv_data <=  -44;
			when -692 => sin_inv_data <=  -44;
			when -691 => sin_inv_data <=  -44;
			when -690 => sin_inv_data <=  -44;
			when -689 => sin_inv_data <=  -44;
			when -688 => sin_inv_data <=  -43;
			when -687 => sin_inv_data <=  -43;
			when -686 => sin_inv_data <=  -43;
			when -685 => sin_inv_data <=  -43;
			when -684 => sin_inv_data <=  -43;
			when -683 => sin_inv_data <=  -43;
			when -682 => sin_inv_data <=  -43;
			when -681 => sin_inv_data <=  -43;
			when -680 => sin_inv_data <=  -43;
			when -679 => sin_inv_data <=  -43;
			when -678 => sin_inv_data <=  -43;
			when -677 => sin_inv_data <=  -43;
			when -676 => sin_inv_data <=  -43;
			when -675 => sin_inv_data <=  -42;
			when -674 => sin_inv_data <=  -42;
			when -673 => sin_inv_data <=  -42;
			when -672 => sin_inv_data <=  -42;
			when -671 => sin_inv_data <=  -42;
			when -670 => sin_inv_data <=  -42;
			when -669 => sin_inv_data <=  -42;
			when -668 => sin_inv_data <=  -42;
			when -667 => sin_inv_data <=  -42;
			when -666 => sin_inv_data <=  -42;
			when -665 => sin_inv_data <=  -42;
			when -664 => sin_inv_data <=  -42;
			when -663 => sin_inv_data <=  -42;
			when -662 => sin_inv_data <=  -41;
			when -661 => sin_inv_data <=  -41;
			when -660 => sin_inv_data <=  -41;
			when -659 => sin_inv_data <=  -41;
			when -658 => sin_inv_data <=  -41;
			when -657 => sin_inv_data <=  -41;
			when -656 => sin_inv_data <=  -41;
			when -655 => sin_inv_data <=  -41;
			when -654 => sin_inv_data <=  -41;
			when -653 => sin_inv_data <=  -41;
			when -652 => sin_inv_data <=  -41;
			when -651 => sin_inv_data <=  -41;
			when -650 => sin_inv_data <=  -41;
			when -649 => sin_inv_data <=  -40;
			when -648 => sin_inv_data <=  -40;
			when -647 => sin_inv_data <=  -40;
			when -646 => sin_inv_data <=  -40;
			when -645 => sin_inv_data <=  -40;
			when -644 => sin_inv_data <=  -40;
			when -643 => sin_inv_data <=  -40;
			when -642 => sin_inv_data <=  -40;
			when -641 => sin_inv_data <=  -40;
			when -640 => sin_inv_data <=  -40;
			when -639 => sin_inv_data <=  -40;
			when -638 => sin_inv_data <=  -40;
			when -637 => sin_inv_data <=  -40;
			when -636 => sin_inv_data <=  -39;
			when -635 => sin_inv_data <=  -39;
			when -634 => sin_inv_data <=  -39;
			when -633 => sin_inv_data <=  -39;
			when -632 => sin_inv_data <=  -39;
			when -631 => sin_inv_data <=  -39;
			when -630 => sin_inv_data <=  -39;
			when -629 => sin_inv_data <=  -39;
			when -628 => sin_inv_data <=  -39;
			when -627 => sin_inv_data <=  -39;
			when -626 => sin_inv_data <=  -39;
			when -625 => sin_inv_data <=  -39;
			when -624 => sin_inv_data <=  -39;
			when -623 => sin_inv_data <=  -39;
			when -622 => sin_inv_data <=  -38;
			when -621 => sin_inv_data <=  -38;
			when -620 => sin_inv_data <=  -38;
			when -619 => sin_inv_data <=  -38;
			when -618 => sin_inv_data <=  -38;
			when -617 => sin_inv_data <=  -38;
			when -616 => sin_inv_data <=  -38;
			when -615 => sin_inv_data <=  -38;
			when -614 => sin_inv_data <=  -38;
			when -613 => sin_inv_data <=  -38;
			when -612 => sin_inv_data <=  -38;
			when -611 => sin_inv_data <=  -38;
			when -610 => sin_inv_data <=  -38;
			when -609 => sin_inv_data <=  -38;
			when -608 => sin_inv_data <=  -37;
			when -607 => sin_inv_data <=  -37;
			when -606 => sin_inv_data <=  -37;
			when -605 => sin_inv_data <=  -37;
			when -604 => sin_inv_data <=  -37;
			when -603 => sin_inv_data <=  -37;
			when -602 => sin_inv_data <=  -37;
			when -601 => sin_inv_data <=  -37;
			when -600 => sin_inv_data <=  -37;
			when -599 => sin_inv_data <=  -37;
			when -598 => sin_inv_data <=  -37;
			when -597 => sin_inv_data <=  -37;
			when -596 => sin_inv_data <=  -37;
			when -595 => sin_inv_data <=  -37;
			when -594 => sin_inv_data <=  -36;
			when -593 => sin_inv_data <=  -36;
			when -592 => sin_inv_data <=  -36;
			when -591 => sin_inv_data <=  -36;
			when -590 => sin_inv_data <=  -36;
			when -589 => sin_inv_data <=  -36;
			when -588 => sin_inv_data <=  -36;
			when -587 => sin_inv_data <=  -36;
			when -586 => sin_inv_data <=  -36;
			when -585 => sin_inv_data <=  -36;
			when -584 => sin_inv_data <=  -36;
			when -583 => sin_inv_data <=  -36;
			when -582 => sin_inv_data <=  -36;
			when -581 => sin_inv_data <=  -36;
			when -580 => sin_inv_data <=  -35;
			when -579 => sin_inv_data <=  -35;
			when -578 => sin_inv_data <=  -35;
			when -577 => sin_inv_data <=  -35;
			when -576 => sin_inv_data <=  -35;
			when -575 => sin_inv_data <=  -35;
			when -574 => sin_inv_data <=  -35;
			when -573 => sin_inv_data <=  -35;
			when -572 => sin_inv_data <=  -35;
			when -571 => sin_inv_data <=  -35;
			when -570 => sin_inv_data <=  -35;
			when -569 => sin_inv_data <=  -35;
			when -568 => sin_inv_data <=  -35;
			when -567 => sin_inv_data <=  -35;
			when -566 => sin_inv_data <=  -34;
			when -565 => sin_inv_data <=  -34;
			when -564 => sin_inv_data <=  -34;
			when -563 => sin_inv_data <=  -34;
			when -562 => sin_inv_data <=  -34;
			when -561 => sin_inv_data <=  -34;
			when -560 => sin_inv_data <=  -34;
			when -559 => sin_inv_data <=  -34;
			when -558 => sin_inv_data <=  -34;
			when -557 => sin_inv_data <=  -34;
			when -556 => sin_inv_data <=  -34;
			when -555 => sin_inv_data <=  -34;
			when -554 => sin_inv_data <=  -34;
			when -553 => sin_inv_data <=  -34;
			when -552 => sin_inv_data <=  -34;
			when -551 => sin_inv_data <=  -33;
			when -550 => sin_inv_data <=  -33;
			when -549 => sin_inv_data <=  -33;
			when -548 => sin_inv_data <=  -33;
			when -547 => sin_inv_data <=  -33;
			when -546 => sin_inv_data <=  -33;
			when -545 => sin_inv_data <=  -33;
			when -544 => sin_inv_data <=  -33;
			when -543 => sin_inv_data <=  -33;
			when -542 => sin_inv_data <=  -33;
			when -541 => sin_inv_data <=  -33;
			when -540 => sin_inv_data <=  -33;
			when -539 => sin_inv_data <=  -33;
			when -538 => sin_inv_data <=  -33;
			when -537 => sin_inv_data <=  -32;
			when -536 => sin_inv_data <=  -32;
			when -535 => sin_inv_data <=  -32;
			when -534 => sin_inv_data <=  -32;
			when -533 => sin_inv_data <=  -32;
			when -532 => sin_inv_data <=  -32;
			when -531 => sin_inv_data <=  -32;
			when -530 => sin_inv_data <=  -32;
			when -529 => sin_inv_data <=  -32;
			when -528 => sin_inv_data <=  -32;
			when -527 => sin_inv_data <=  -32;
			when -526 => sin_inv_data <=  -32;
			when -525 => sin_inv_data <=  -32;
			when -524 => sin_inv_data <=  -32;
			when -523 => sin_inv_data <=  -32;
			when -522 => sin_inv_data <=  -31;
			when -521 => sin_inv_data <=  -31;
			when -520 => sin_inv_data <=  -31;
			when -519 => sin_inv_data <=  -31;
			when -518 => sin_inv_data <=  -31;
			when -517 => sin_inv_data <=  -31;
			when -516 => sin_inv_data <=  -31;
			when -515 => sin_inv_data <=  -31;
			when -514 => sin_inv_data <=  -31;
			when -513 => sin_inv_data <=  -31;
			when -512 => sin_inv_data <=  -31;
			when -511 => sin_inv_data <=  -31;
			when -510 => sin_inv_data <=  -31;
			when -509 => sin_inv_data <=  -31;
			when -508 => sin_inv_data <=  -31;
			when -507 => sin_inv_data <=  -30;
			when -506 => sin_inv_data <=  -30;
			when -505 => sin_inv_data <=  -30;
			when -504 => sin_inv_data <=  -30;
			when -503 => sin_inv_data <=  -30;
			when -502 => sin_inv_data <=  -30;
			when -501 => sin_inv_data <=  -30;
			when -500 => sin_inv_data <=  -30;
			when -499 => sin_inv_data <=  -30;
			when -498 => sin_inv_data <=  -30;
			when -497 => sin_inv_data <=  -30;
			when -496 => sin_inv_data <=  -30;
			when -495 => sin_inv_data <=  -30;
			when -494 => sin_inv_data <=  -30;
			when -493 => sin_inv_data <=  -30;
			when -492 => sin_inv_data <=  -29;
			when -491 => sin_inv_data <=  -29;
			when -490 => sin_inv_data <=  -29;
			when -489 => sin_inv_data <=  -29;
			when -488 => sin_inv_data <=  -29;
			when -487 => sin_inv_data <=  -29;
			when -486 => sin_inv_data <=  -29;
			when -485 => sin_inv_data <=  -29;
			when -484 => sin_inv_data <=  -29;
			when -483 => sin_inv_data <=  -29;
			when -482 => sin_inv_data <=  -29;
			when -481 => sin_inv_data <=  -29;
			when -480 => sin_inv_data <=  -29;
			when -479 => sin_inv_data <=  -29;
			when -478 => sin_inv_data <=  -29;
			when -477 => sin_inv_data <=  -28;
			when -476 => sin_inv_data <=  -28;
			when -475 => sin_inv_data <=  -28;
			when -474 => sin_inv_data <=  -28;
			when -473 => sin_inv_data <=  -28;
			when -472 => sin_inv_data <=  -28;
			when -471 => sin_inv_data <=  -28;
			when -470 => sin_inv_data <=  -28;
			when -469 => sin_inv_data <=  -28;
			when -468 => sin_inv_data <=  -28;
			when -467 => sin_inv_data <=  -28;
			when -466 => sin_inv_data <=  -28;
			when -465 => sin_inv_data <=  -28;
			when -464 => sin_inv_data <=  -28;
			when -463 => sin_inv_data <=  -28;
			when -462 => sin_inv_data <=  -28;
			when -461 => sin_inv_data <=  -27;
			when -460 => sin_inv_data <=  -27;
			when -459 => sin_inv_data <=  -27;
			when -458 => sin_inv_data <=  -27;
			when -457 => sin_inv_data <=  -27;
			when -456 => sin_inv_data <=  -27;
			when -455 => sin_inv_data <=  -27;
			when -454 => sin_inv_data <=  -27;
			when -453 => sin_inv_data <=  -27;
			when -452 => sin_inv_data <=  -27;
			when -451 => sin_inv_data <=  -27;
			when -450 => sin_inv_data <=  -27;
			when -449 => sin_inv_data <=  -27;
			when -448 => sin_inv_data <=  -27;
			when -447 => sin_inv_data <=  -27;
			when -446 => sin_inv_data <=  -26;
			when -445 => sin_inv_data <=  -26;
			when -444 => sin_inv_data <=  -26;
			when -443 => sin_inv_data <=  -26;
			when -442 => sin_inv_data <=  -26;
			when -441 => sin_inv_data <=  -26;
			when -440 => sin_inv_data <=  -26;
			when -439 => sin_inv_data <=  -26;
			when -438 => sin_inv_data <=  -26;
			when -437 => sin_inv_data <=  -26;
			when -436 => sin_inv_data <=  -26;
			when -435 => sin_inv_data <=  -26;
			when -434 => sin_inv_data <=  -26;
			when -433 => sin_inv_data <=  -26;
			when -432 => sin_inv_data <=  -26;
			when -431 => sin_inv_data <=  -26;
			when -430 => sin_inv_data <=  -25;
			when -429 => sin_inv_data <=  -25;
			when -428 => sin_inv_data <=  -25;
			when -427 => sin_inv_data <=  -25;
			when -426 => sin_inv_data <=  -25;
			when -425 => sin_inv_data <=  -25;
			when -424 => sin_inv_data <=  -25;
			when -423 => sin_inv_data <=  -25;
			when -422 => sin_inv_data <=  -25;
			when -421 => sin_inv_data <=  -25;
			when -420 => sin_inv_data <=  -25;
			when -419 => sin_inv_data <=  -25;
			when -418 => sin_inv_data <=  -25;
			when -417 => sin_inv_data <=  -25;
			when -416 => sin_inv_data <=  -25;
			when -415 => sin_inv_data <=  -25;
			when -414 => sin_inv_data <=  -24;
			when -413 => sin_inv_data <=  -24;
			when -412 => sin_inv_data <=  -24;
			when -411 => sin_inv_data <=  -24;
			when -410 => sin_inv_data <=  -24;
			when -409 => sin_inv_data <=  -24;
			when -408 => sin_inv_data <=  -24;
			when -407 => sin_inv_data <=  -24;
			when -406 => sin_inv_data <=  -24;
			when -405 => sin_inv_data <=  -24;
			when -404 => sin_inv_data <=  -24;
			when -403 => sin_inv_data <=  -24;
			when -402 => sin_inv_data <=  -24;
			when -401 => sin_inv_data <=  -24;
			when -400 => sin_inv_data <=  -24;
			when -399 => sin_inv_data <=  -24;
			when -398 => sin_inv_data <=  -23;
			when -397 => sin_inv_data <=  -23;
			when -396 => sin_inv_data <=  -23;
			when -395 => sin_inv_data <=  -23;
			when -394 => sin_inv_data <=  -23;
			when -393 => sin_inv_data <=  -23;
			when -392 => sin_inv_data <=  -23;
			when -391 => sin_inv_data <=  -23;
			when -390 => sin_inv_data <=  -23;
			when -389 => sin_inv_data <=  -23;
			when -388 => sin_inv_data <=  -23;
			when -387 => sin_inv_data <=  -23;
			when -386 => sin_inv_data <=  -23;
			when -385 => sin_inv_data <=  -23;
			when -384 => sin_inv_data <=  -23;
			when -383 => sin_inv_data <=  -23;
			when -382 => sin_inv_data <=  -22;
			when -381 => sin_inv_data <=  -22;
			when -380 => sin_inv_data <=  -22;
			when -379 => sin_inv_data <=  -22;
			when -378 => sin_inv_data <=  -22;
			when -377 => sin_inv_data <=  -22;
			when -376 => sin_inv_data <=  -22;
			when -375 => sin_inv_data <=  -22;
			when -374 => sin_inv_data <=  -22;
			when -373 => sin_inv_data <=  -22;
			when -372 => sin_inv_data <=  -22;
			when -371 => sin_inv_data <=  -22;
			when -370 => sin_inv_data <=  -22;
			when -369 => sin_inv_data <=  -22;
			when -368 => sin_inv_data <=  -22;
			when -367 => sin_inv_data <=  -22;
			when -366 => sin_inv_data <=  -21;
			when -365 => sin_inv_data <=  -21;
			when -364 => sin_inv_data <=  -21;
			when -363 => sin_inv_data <=  -21;
			when -362 => sin_inv_data <=  -21;
			when -361 => sin_inv_data <=  -21;
			when -360 => sin_inv_data <=  -21;
			when -359 => sin_inv_data <=  -21;
			when -358 => sin_inv_data <=  -21;
			when -357 => sin_inv_data <=  -21;
			when -356 => sin_inv_data <=  -21;
			when -355 => sin_inv_data <=  -21;
			when -354 => sin_inv_data <=  -21;
			when -353 => sin_inv_data <=  -21;
			when -352 => sin_inv_data <=  -21;
			when -351 => sin_inv_data <=  -21;
			when -350 => sin_inv_data <=  -20;
			when -349 => sin_inv_data <=  -20;
			when -348 => sin_inv_data <=  -20;
			when -347 => sin_inv_data <=  -20;
			when -346 => sin_inv_data <=  -20;
			when -345 => sin_inv_data <=  -20;
			when -344 => sin_inv_data <=  -20;
			when -343 => sin_inv_data <=  -20;
			when -342 => sin_inv_data <=  -20;
			when -341 => sin_inv_data <=  -20;
			when -340 => sin_inv_data <=  -20;
			when -339 => sin_inv_data <=  -20;
			when -338 => sin_inv_data <=  -20;
			when -337 => sin_inv_data <=  -20;
			when -336 => sin_inv_data <=  -20;
			when -335 => sin_inv_data <=  -20;
			when -334 => sin_inv_data <=  -20;
			when -333 => sin_inv_data <=  -19;
			when -332 => sin_inv_data <=  -19;
			when -331 => sin_inv_data <=  -19;
			when -330 => sin_inv_data <=  -19;
			when -329 => sin_inv_data <=  -19;
			when -328 => sin_inv_data <=  -19;
			when -327 => sin_inv_data <=  -19;
			when -326 => sin_inv_data <=  -19;
			when -325 => sin_inv_data <=  -19;
			when -324 => sin_inv_data <=  -19;
			when -323 => sin_inv_data <=  -19;
			when -322 => sin_inv_data <=  -19;
			when -321 => sin_inv_data <=  -19;
			when -320 => sin_inv_data <=  -19;
			when -319 => sin_inv_data <=  -19;
			when -318 => sin_inv_data <=  -19;
			when -317 => sin_inv_data <=  -18;
			when -316 => sin_inv_data <=  -18;
			when -315 => sin_inv_data <=  -18;
			when -314 => sin_inv_data <=  -18;
			when -313 => sin_inv_data <=  -18;
			when -312 => sin_inv_data <=  -18;
			when -311 => sin_inv_data <=  -18;
			when -310 => sin_inv_data <=  -18;
			when -309 => sin_inv_data <=  -18;
			when -308 => sin_inv_data <=  -18;
			when -307 => sin_inv_data <=  -18;
			when -306 => sin_inv_data <=  -18;
			when -305 => sin_inv_data <=  -18;
			when -304 => sin_inv_data <=  -18;
			when -303 => sin_inv_data <=  -18;
			when -302 => sin_inv_data <=  -18;
			when -301 => sin_inv_data <=  -18;
			when -300 => sin_inv_data <=  -17;
			when -299 => sin_inv_data <=  -17;
			when -298 => sin_inv_data <=  -17;
			when -297 => sin_inv_data <=  -17;
			when -296 => sin_inv_data <=  -17;
			when -295 => sin_inv_data <=  -17;
			when -294 => sin_inv_data <=  -17;
			when -293 => sin_inv_data <=  -17;
			when -292 => sin_inv_data <=  -17;
			when -291 => sin_inv_data <=  -17;
			when -290 => sin_inv_data <=  -17;
			when -289 => sin_inv_data <=  -17;
			when -288 => sin_inv_data <=  -17;
			when -287 => sin_inv_data <=  -17;
			when -286 => sin_inv_data <=  -17;
			when -285 => sin_inv_data <=  -17;
			when -284 => sin_inv_data <=  -16;
			when -283 => sin_inv_data <=  -16;
			when -282 => sin_inv_data <=  -16;
			when -281 => sin_inv_data <=  -16;
			when -280 => sin_inv_data <=  -16;
			when -279 => sin_inv_data <=  -16;
			when -278 => sin_inv_data <=  -16;
			when -277 => sin_inv_data <=  -16;
			when -276 => sin_inv_data <=  -16;
			when -275 => sin_inv_data <=  -16;
			when -274 => sin_inv_data <=  -16;
			when -273 => sin_inv_data <=  -16;
			when -272 => sin_inv_data <=  -16;
			when -271 => sin_inv_data <=  -16;
			when -270 => sin_inv_data <=  -16;
			when -269 => sin_inv_data <=  -16;
			when -268 => sin_inv_data <=  -16;
			when -267 => sin_inv_data <=  -15;
			when -266 => sin_inv_data <=  -15;
			when -265 => sin_inv_data <=  -15;
			when -264 => sin_inv_data <=  -15;
			when -263 => sin_inv_data <=  -15;
			when -262 => sin_inv_data <=  -15;
			when -261 => sin_inv_data <=  -15;
			when -260 => sin_inv_data <=  -15;
			when -259 => sin_inv_data <=  -15;
			when -258 => sin_inv_data <=  -15;
			when -257 => sin_inv_data <=  -15;
			when -256 => sin_inv_data <=  -15;
			when -255 => sin_inv_data <=  -15;
			when -254 => sin_inv_data <=  -15;
			when -253 => sin_inv_data <=  -15;
			when -252 => sin_inv_data <=  -15;
			when -251 => sin_inv_data <=  -15;
			when -250 => sin_inv_data <=  -14;
			when -249 => sin_inv_data <=  -14;
			when -248 => sin_inv_data <=  -14;
			when -247 => sin_inv_data <=  -14;
			when -246 => sin_inv_data <=  -14;
			when -245 => sin_inv_data <=  -14;
			when -244 => sin_inv_data <=  -14;
			when -243 => sin_inv_data <=  -14;
			when -242 => sin_inv_data <=  -14;
			when -241 => sin_inv_data <=  -14;
			when -240 => sin_inv_data <=  -14;
			when -239 => sin_inv_data <=  -14;
			when -238 => sin_inv_data <=  -14;
			when -237 => sin_inv_data <=  -14;
			when -236 => sin_inv_data <=  -14;
			when -235 => sin_inv_data <=  -14;
			when -234 => sin_inv_data <=  -14;
			when -233 => sin_inv_data <=  -13;
			when -232 => sin_inv_data <=  -13;
			when -231 => sin_inv_data <=  -13;
			when -230 => sin_inv_data <=  -13;
			when -229 => sin_inv_data <=  -13;
			when -228 => sin_inv_data <=  -13;
			when -227 => sin_inv_data <=  -13;
			when -226 => sin_inv_data <=  -13;
			when -225 => sin_inv_data <=  -13;
			when -224 => sin_inv_data <=  -13;
			when -223 => sin_inv_data <=  -13;
			when -222 => sin_inv_data <=  -13;
			when -221 => sin_inv_data <=  -13;
			when -220 => sin_inv_data <=  -13;
			when -219 => sin_inv_data <=  -13;
			when -218 => sin_inv_data <=  -13;
			when -217 => sin_inv_data <=  -13;
			when -216 => sin_inv_data <=  -12;
			when -215 => sin_inv_data <=  -12;
			when -214 => sin_inv_data <=  -12;
			when -213 => sin_inv_data <=  -12;
			when -212 => sin_inv_data <=  -12;
			when -211 => sin_inv_data <=  -12;
			when -210 => sin_inv_data <=  -12;
			when -209 => sin_inv_data <=  -12;
			when -208 => sin_inv_data <=  -12;
			when -207 => sin_inv_data <=  -12;
			when -206 => sin_inv_data <=  -12;
			when -205 => sin_inv_data <=  -12;
			when -204 => sin_inv_data <=  -12;
			when -203 => sin_inv_data <=  -12;
			when -202 => sin_inv_data <=  -12;
			when -201 => sin_inv_data <=  -12;
			when -200 => sin_inv_data <=  -12;
			when -199 => sin_inv_data <=  -11;
			when -198 => sin_inv_data <=  -11;
			when -197 => sin_inv_data <=  -11;
			when -196 => sin_inv_data <=  -11;
			when -195 => sin_inv_data <=  -11;
			when -194 => sin_inv_data <=  -11;
			when -193 => sin_inv_data <=  -11;
			when -192 => sin_inv_data <=  -11;
			when -191 => sin_inv_data <=  -11;
			when -190 => sin_inv_data <=  -11;
			when -189 => sin_inv_data <=  -11;
			when -188 => sin_inv_data <=  -11;
			when -187 => sin_inv_data <=  -11;
			when -186 => sin_inv_data <=  -11;
			when -185 => sin_inv_data <=  -11;
			when -184 => sin_inv_data <=  -11;
			when -183 => sin_inv_data <=  -11;
			when -182 => sin_inv_data <=  -10;
			when -181 => sin_inv_data <=  -10;
			when -180 => sin_inv_data <=  -10;
			when -179 => sin_inv_data <=  -10;
			when -178 => sin_inv_data <=  -10;
			when -177 => sin_inv_data <=  -10;
			when -176 => sin_inv_data <=  -10;
			when -175 => sin_inv_data <=  -10;
			when -174 => sin_inv_data <=  -10;
			when -173 => sin_inv_data <=  -10;
			when -172 => sin_inv_data <=  -10;
			when -171 => sin_inv_data <=  -10;
			when -170 => sin_inv_data <=  -10;
			when -169 => sin_inv_data <=  -10;
			when -168 => sin_inv_data <=  -10;
			when -167 => sin_inv_data <=  -10;
			when -166 => sin_inv_data <=  -10;
			when -165 => sin_inv_data <=  -9;
			when -164 => sin_inv_data <=  -9;
			when -163 => sin_inv_data <=  -9;
			when -162 => sin_inv_data <=  -9;
			when -161 => sin_inv_data <=  -9;
			when -160 => sin_inv_data <=  -9;
			when -159 => sin_inv_data <=  -9;
			when -158 => sin_inv_data <=  -9;
			when -157 => sin_inv_data <=  -9;
			when -156 => sin_inv_data <=  -9;
			when -155 => sin_inv_data <=  -9;
			when -154 => sin_inv_data <=  -9;
			when -153 => sin_inv_data <=  -9;
			when -152 => sin_inv_data <=  -9;
			when -151 => sin_inv_data <=  -9;
			when -150 => sin_inv_data <=  -9;
			when -149 => sin_inv_data <=  -9;
			when -148 => sin_inv_data <=  -9;
			when -147 => sin_inv_data <=  -8;
			when -146 => sin_inv_data <=  -8;
			when -145 => sin_inv_data <=  -8;
			when -144 => sin_inv_data <=  -8;
			when -143 => sin_inv_data <=  -8;
			when -142 => sin_inv_data <=  -8;
			when -141 => sin_inv_data <=  -8;
			when -140 => sin_inv_data <=  -8;
			when -139 => sin_inv_data <=  -8;
			when -138 => sin_inv_data <=  -8;
			when -137 => sin_inv_data <=  -8;
			when -136 => sin_inv_data <=  -8;
			when -135 => sin_inv_data <=  -8;
			when -134 => sin_inv_data <=  -8;
			when -133 => sin_inv_data <=  -8;
			when -132 => sin_inv_data <=  -8;
			when -131 => sin_inv_data <=  -8;
			when -130 => sin_inv_data <=  -7;
			when -129 => sin_inv_data <=  -7;
			when -128 => sin_inv_data <=  -7;
			when -127 => sin_inv_data <=  -7;
			when -126 => sin_inv_data <=  -7;
			when -125 => sin_inv_data <=  -7;
			when -124 => sin_inv_data <=  -7;
			when -123 => sin_inv_data <=  -7;
			when -122 => sin_inv_data <=  -7;
			when -121 => sin_inv_data <=  -7;
			when -120 => sin_inv_data <=  -7;
			when -119 => sin_inv_data <=  -7;
			when -118 => sin_inv_data <=  -7;
			when -117 => sin_inv_data <=  -7;
			when -116 => sin_inv_data <=  -7;
			when -115 => sin_inv_data <=  -7;
			when -114 => sin_inv_data <=  -7;
			when -113 => sin_inv_data <=  -6;
			when -112 => sin_inv_data <=  -6;
			when -111 => sin_inv_data <=  -6;
			when -110 => sin_inv_data <=  -6;
			when -109 => sin_inv_data <=  -6;
			when -108 => sin_inv_data <=  -6;
			when -107 => sin_inv_data <=  -6;
			when -106 => sin_inv_data <=  -6;
			when -105 => sin_inv_data <=  -6;
			when -104 => sin_inv_data <=  -6;
			when -103 => sin_inv_data <=  -6;
			when -102 => sin_inv_data <=  -6;
			when -101 => sin_inv_data <=  -6;
			when -100 => sin_inv_data <=  -6;
			when -99 => sin_inv_data <=  -6;
			when -98 => sin_inv_data <=  -6;
			when -97 => sin_inv_data <=  -6;
			when -96 => sin_inv_data <=  -6;
			when -95 => sin_inv_data <=  -5;
			when -94 => sin_inv_data <=  -5;
			when -93 => sin_inv_data <=  -5;
			when -92 => sin_inv_data <=  -5;
			when -91 => sin_inv_data <=  -5;
			when -90 => sin_inv_data <=  -5;
			when -89 => sin_inv_data <=  -5;
			when -88 => sin_inv_data <=  -5;
			when -87 => sin_inv_data <=  -5;
			when -86 => sin_inv_data <=  -5;
			when -85 => sin_inv_data <=  -5;
			when -84 => sin_inv_data <=  -5;
			when -83 => sin_inv_data <=  -5;
			when -82 => sin_inv_data <=  -5;
			when -81 => sin_inv_data <=  -5;
			when -80 => sin_inv_data <=  -5;
			when -79 => sin_inv_data <=  -5;
			when -78 => sin_inv_data <=  -4;
			when -77 => sin_inv_data <=  -4;
			when -76 => sin_inv_data <=  -4;
			when -75 => sin_inv_data <=  -4;
			when -74 => sin_inv_data <=  -4;
			when -73 => sin_inv_data <=  -4;
			when -72 => sin_inv_data <=  -4;
			when -71 => sin_inv_data <=  -4;
			when -70 => sin_inv_data <=  -4;
			when -69 => sin_inv_data <=  -4;
			when -68 => sin_inv_data <=  -4;
			when -67 => sin_inv_data <=  -4;
			when -66 => sin_inv_data <=  -4;
			when -65 => sin_inv_data <=  -4;
			when -64 => sin_inv_data <=  -4;
			when -63 => sin_inv_data <=  -4;
			when -62 => sin_inv_data <=  -4;
			when -61 => sin_inv_data <=  -3;
			when -60 => sin_inv_data <=  -3;
			when -59 => sin_inv_data <=  -3;
			when -58 => sin_inv_data <=  -3;
			when -57 => sin_inv_data <=  -3;
			when -56 => sin_inv_data <=  -3;
			when -55 => sin_inv_data <=  -3;
			when -54 => sin_inv_data <=  -3;
			when -53 => sin_inv_data <=  -3;
			when -52 => sin_inv_data <=  -3;
			when -51 => sin_inv_data <=  -3;
			when -50 => sin_inv_data <=  -3;
			when -49 => sin_inv_data <=  -3;
			when -48 => sin_inv_data <=  -3;
			when -47 => sin_inv_data <=  -3;
			when -46 => sin_inv_data <=  -3;
			when -45 => sin_inv_data <=  -3;
			when -44 => sin_inv_data <=  -3;
			when -43 => sin_inv_data <=  -2;
			when -42 => sin_inv_data <=  -2;
			when -41 => sin_inv_data <=  -2;
			when -40 => sin_inv_data <=  -2;
			when -39 => sin_inv_data <=  -2;
			when -38 => sin_inv_data <=  -2;
			when -37 => sin_inv_data <=  -2;
			when -36 => sin_inv_data <=  -2;
			when -35 => sin_inv_data <=  -2;
			when -34 => sin_inv_data <=  -2;
			when -33 => sin_inv_data <=  -2;
			when -32 => sin_inv_data <=  -2;
			when -31 => sin_inv_data <=  -2;
			when -30 => sin_inv_data <=  -2;
			when -29 => sin_inv_data <=  -2;
			when -28 => sin_inv_data <=  -2;
			when -27 => sin_inv_data <=  -2;
			when -26 => sin_inv_data <=  -1;
			when -25 => sin_inv_data <=  -1;
			when -24 => sin_inv_data <=  -1;
			when -23 => sin_inv_data <=  -1;
			when -22 => sin_inv_data <=  -1;
			when -21 => sin_inv_data <=  -1;
			when -20 => sin_inv_data <=  -1;
			when -19 => sin_inv_data <=  -1;
			when -18 => sin_inv_data <=  -1;
			when -17 => sin_inv_data <=  -1;
			when -16 => sin_inv_data <=  -1;
			when -15 => sin_inv_data <=  -1;
			when -14 => sin_inv_data <=  -1;
			when -13 => sin_inv_data <=  -1;
			when -12 => sin_inv_data <=  -1;
			when -11 => sin_inv_data <=  -1;
			when -10 => sin_inv_data <=  -1;
			when -9 => sin_inv_data <=  -1;
			when -8 => sin_inv_data <=  0;
			when -7 => sin_inv_data <=  0;
			when -6 => sin_inv_data <=  0;
			when -5 => sin_inv_data <=  0;
			when -4 => sin_inv_data <=  0;
			when -3 => sin_inv_data <=  0;
			when -2 => sin_inv_data <=  0;
			when -1 => sin_inv_data <=  0;
			when 0 => sin_inv_data <=  0;
			when 1 => sin_inv_data <=  0;
			when 2 => sin_inv_data <=  0;
			when 3 => sin_inv_data <=  0;
			when 4 => sin_inv_data <=  0;
			when 5 => sin_inv_data <=  0;
			when 6 => sin_inv_data <=  0;
			when 7 => sin_inv_data <=  0;
			when 8 => sin_inv_data <=  0;
			when 9 => sin_inv_data <=  1;
			when 10 => sin_inv_data <=  1;
			when 11 => sin_inv_data <=  1;
			when 12 => sin_inv_data <=  1;
			when 13 => sin_inv_data <=  1;
			when 14 => sin_inv_data <=  1;
			when 15 => sin_inv_data <=  1;
			when 16 => sin_inv_data <=  1;
			when 17 => sin_inv_data <=  1;
			when 18 => sin_inv_data <=  1;
			when 19 => sin_inv_data <=  1;
			when 20 => sin_inv_data <=  1;
			when 21 => sin_inv_data <=  1;
			when 22 => sin_inv_data <=  1;
			when 23 => sin_inv_data <=  1;
			when 24 => sin_inv_data <=  1;
			when 25 => sin_inv_data <=  1;
			when 26 => sin_inv_data <=  1;
			when 27 => sin_inv_data <=  2;
			when 28 => sin_inv_data <=  2;
			when 29 => sin_inv_data <=  2;
			when 30 => sin_inv_data <=  2;
			when 31 => sin_inv_data <=  2;
			when 32 => sin_inv_data <=  2;
			when 33 => sin_inv_data <=  2;
			when 34 => sin_inv_data <=  2;
			when 35 => sin_inv_data <=  2;
			when 36 => sin_inv_data <=  2;
			when 37 => sin_inv_data <=  2;
			when 38 => sin_inv_data <=  2;
			when 39 => sin_inv_data <=  2;
			when 40 => sin_inv_data <=  2;
			when 41 => sin_inv_data <=  2;
			when 42 => sin_inv_data <=  2;
			when 43 => sin_inv_data <=  2;
			when 44 => sin_inv_data <=  3;
			when 45 => sin_inv_data <=  3;
			when 46 => sin_inv_data <=  3;
			when 47 => sin_inv_data <=  3;
			when 48 => sin_inv_data <=  3;
			when 49 => sin_inv_data <=  3;
			when 50 => sin_inv_data <=  3;
			when 51 => sin_inv_data <=  3;
			when 52 => sin_inv_data <=  3;
			when 53 => sin_inv_data <=  3;
			when 54 => sin_inv_data <=  3;
			when 55 => sin_inv_data <=  3;
			when 56 => sin_inv_data <=  3;
			when 57 => sin_inv_data <=  3;
			when 58 => sin_inv_data <=  3;
			when 59 => sin_inv_data <=  3;
			when 60 => sin_inv_data <=  3;
			when 61 => sin_inv_data <=  3;
			when 62 => sin_inv_data <=  4;
			when 63 => sin_inv_data <=  4;
			when 64 => sin_inv_data <=  4;
			when 65 => sin_inv_data <=  4;
			when 66 => sin_inv_data <=  4;
			when 67 => sin_inv_data <=  4;
			when 68 => sin_inv_data <=  4;
			when 69 => sin_inv_data <=  4;
			when 70 => sin_inv_data <=  4;
			when 71 => sin_inv_data <=  4;
			when 72 => sin_inv_data <=  4;
			when 73 => sin_inv_data <=  4;
			when 74 => sin_inv_data <=  4;
			when 75 => sin_inv_data <=  4;
			when 76 => sin_inv_data <=  4;
			when 77 => sin_inv_data <=  4;
			when 78 => sin_inv_data <=  4;
			when 79 => sin_inv_data <=  5;
			when 80 => sin_inv_data <=  5;
			when 81 => sin_inv_data <=  5;
			when 82 => sin_inv_data <=  5;
			when 83 => sin_inv_data <=  5;
			when 84 => sin_inv_data <=  5;
			when 85 => sin_inv_data <=  5;
			when 86 => sin_inv_data <=  5;
			when 87 => sin_inv_data <=  5;
			when 88 => sin_inv_data <=  5;
			when 89 => sin_inv_data <=  5;
			when 90 => sin_inv_data <=  5;
			when 91 => sin_inv_data <=  5;
			when 92 => sin_inv_data <=  5;
			when 93 => sin_inv_data <=  5;
			when 94 => sin_inv_data <=  5;
			when 95 => sin_inv_data <=  5;
			when 96 => sin_inv_data <=  6;
			when 97 => sin_inv_data <=  6;
			when 98 => sin_inv_data <=  6;
			when 99 => sin_inv_data <=  6;
			when 100 => sin_inv_data <=  6;
			when 101 => sin_inv_data <=  6;
			when 102 => sin_inv_data <=  6;
			when 103 => sin_inv_data <=  6;
			when 104 => sin_inv_data <=  6;
			when 105 => sin_inv_data <=  6;
			when 106 => sin_inv_data <=  6;
			when 107 => sin_inv_data <=  6;
			when 108 => sin_inv_data <=  6;
			when 109 => sin_inv_data <=  6;
			when 110 => sin_inv_data <=  6;
			when 111 => sin_inv_data <=  6;
			when 112 => sin_inv_data <=  6;
			when 113 => sin_inv_data <=  6;
			when 114 => sin_inv_data <=  7;
			when 115 => sin_inv_data <=  7;
			when 116 => sin_inv_data <=  7;
			when 117 => sin_inv_data <=  7;
			when 118 => sin_inv_data <=  7;
			when 119 => sin_inv_data <=  7;
			when 120 => sin_inv_data <=  7;
			when 121 => sin_inv_data <=  7;
			when 122 => sin_inv_data <=  7;
			when 123 => sin_inv_data <=  7;
			when 124 => sin_inv_data <=  7;
			when 125 => sin_inv_data <=  7;
			when 126 => sin_inv_data <=  7;
			when 127 => sin_inv_data <=  7;
			when 128 => sin_inv_data <=  7;
			when 129 => sin_inv_data <=  7;
			when 130 => sin_inv_data <=  7;
			when 131 => sin_inv_data <=  8;
			when 132 => sin_inv_data <=  8;
			when 133 => sin_inv_data <=  8;
			when 134 => sin_inv_data <=  8;
			when 135 => sin_inv_data <=  8;
			when 136 => sin_inv_data <=  8;
			when 137 => sin_inv_data <=  8;
			when 138 => sin_inv_data <=  8;
			when 139 => sin_inv_data <=  8;
			when 140 => sin_inv_data <=  8;
			when 141 => sin_inv_data <=  8;
			when 142 => sin_inv_data <=  8;
			when 143 => sin_inv_data <=  8;
			when 144 => sin_inv_data <=  8;
			when 145 => sin_inv_data <=  8;
			when 146 => sin_inv_data <=  8;
			when 147 => sin_inv_data <=  8;
			when 148 => sin_inv_data <=  9;
			when 149 => sin_inv_data <=  9;
			when 150 => sin_inv_data <=  9;
			when 151 => sin_inv_data <=  9;
			when 152 => sin_inv_data <=  9;
			when 153 => sin_inv_data <=  9;
			when 154 => sin_inv_data <=  9;
			when 155 => sin_inv_data <=  9;
			when 156 => sin_inv_data <=  9;
			when 157 => sin_inv_data <=  9;
			when 158 => sin_inv_data <=  9;
			when 159 => sin_inv_data <=  9;
			when 160 => sin_inv_data <=  9;
			when 161 => sin_inv_data <=  9;
			when 162 => sin_inv_data <=  9;
			when 163 => sin_inv_data <=  9;
			when 164 => sin_inv_data <=  9;
			when 165 => sin_inv_data <=  9;
			when 166 => sin_inv_data <=  10;
			when 167 => sin_inv_data <=  10;
			when 168 => sin_inv_data <=  10;
			when 169 => sin_inv_data <=  10;
			when 170 => sin_inv_data <=  10;
			when 171 => sin_inv_data <=  10;
			when 172 => sin_inv_data <=  10;
			when 173 => sin_inv_data <=  10;
			when 174 => sin_inv_data <=  10;
			when 175 => sin_inv_data <=  10;
			when 176 => sin_inv_data <=  10;
			when 177 => sin_inv_data <=  10;
			when 178 => sin_inv_data <=  10;
			when 179 => sin_inv_data <=  10;
			when 180 => sin_inv_data <=  10;
			when 181 => sin_inv_data <=  10;
			when 182 => sin_inv_data <=  10;
			when 183 => sin_inv_data <=  11;
			when 184 => sin_inv_data <=  11;
			when 185 => sin_inv_data <=  11;
			when 186 => sin_inv_data <=  11;
			when 187 => sin_inv_data <=  11;
			when 188 => sin_inv_data <=  11;
			when 189 => sin_inv_data <=  11;
			when 190 => sin_inv_data <=  11;
			when 191 => sin_inv_data <=  11;
			when 192 => sin_inv_data <=  11;
			when 193 => sin_inv_data <=  11;
			when 194 => sin_inv_data <=  11;
			when 195 => sin_inv_data <=  11;
			when 196 => sin_inv_data <=  11;
			when 197 => sin_inv_data <=  11;
			when 198 => sin_inv_data <=  11;
			when 199 => sin_inv_data <=  11;
			when 200 => sin_inv_data <=  12;
			when 201 => sin_inv_data <=  12;
			when 202 => sin_inv_data <=  12;
			when 203 => sin_inv_data <=  12;
			when 204 => sin_inv_data <=  12;
			when 205 => sin_inv_data <=  12;
			when 206 => sin_inv_data <=  12;
			when 207 => sin_inv_data <=  12;
			when 208 => sin_inv_data <=  12;
			when 209 => sin_inv_data <=  12;
			when 210 => sin_inv_data <=  12;
			when 211 => sin_inv_data <=  12;
			when 212 => sin_inv_data <=  12;
			when 213 => sin_inv_data <=  12;
			when 214 => sin_inv_data <=  12;
			when 215 => sin_inv_data <=  12;
			when 216 => sin_inv_data <=  12;
			when 217 => sin_inv_data <=  13;
			when 218 => sin_inv_data <=  13;
			when 219 => sin_inv_data <=  13;
			when 220 => sin_inv_data <=  13;
			when 221 => sin_inv_data <=  13;
			when 222 => sin_inv_data <=  13;
			when 223 => sin_inv_data <=  13;
			when 224 => sin_inv_data <=  13;
			when 225 => sin_inv_data <=  13;
			when 226 => sin_inv_data <=  13;
			when 227 => sin_inv_data <=  13;
			when 228 => sin_inv_data <=  13;
			when 229 => sin_inv_data <=  13;
			when 230 => sin_inv_data <=  13;
			when 231 => sin_inv_data <=  13;
			when 232 => sin_inv_data <=  13;
			when 233 => sin_inv_data <=  13;
			when 234 => sin_inv_data <=  14;
			when 235 => sin_inv_data <=  14;
			when 236 => sin_inv_data <=  14;
			when 237 => sin_inv_data <=  14;
			when 238 => sin_inv_data <=  14;
			when 239 => sin_inv_data <=  14;
			when 240 => sin_inv_data <=  14;
			when 241 => sin_inv_data <=  14;
			when 242 => sin_inv_data <=  14;
			when 243 => sin_inv_data <=  14;
			when 244 => sin_inv_data <=  14;
			when 245 => sin_inv_data <=  14;
			when 246 => sin_inv_data <=  14;
			when 247 => sin_inv_data <=  14;
			when 248 => sin_inv_data <=  14;
			when 249 => sin_inv_data <=  14;
			when 250 => sin_inv_data <=  14;
			when 251 => sin_inv_data <=  15;
			when 252 => sin_inv_data <=  15;
			when 253 => sin_inv_data <=  15;
			when 254 => sin_inv_data <=  15;
			when 255 => sin_inv_data <=  15;
			when 256 => sin_inv_data <=  15;
			when 257 => sin_inv_data <=  15;
			when 258 => sin_inv_data <=  15;
			when 259 => sin_inv_data <=  15;
			when 260 => sin_inv_data <=  15;
			when 261 => sin_inv_data <=  15;
			when 262 => sin_inv_data <=  15;
			when 263 => sin_inv_data <=  15;
			when 264 => sin_inv_data <=  15;
			when 265 => sin_inv_data <=  15;
			when 266 => sin_inv_data <=  15;
			when 267 => sin_inv_data <=  15;
			when 268 => sin_inv_data <=  16;
			when 269 => sin_inv_data <=  16;
			when 270 => sin_inv_data <=  16;
			when 271 => sin_inv_data <=  16;
			when 272 => sin_inv_data <=  16;
			when 273 => sin_inv_data <=  16;
			when 274 => sin_inv_data <=  16;
			when 275 => sin_inv_data <=  16;
			when 276 => sin_inv_data <=  16;
			when 277 => sin_inv_data <=  16;
			when 278 => sin_inv_data <=  16;
			when 279 => sin_inv_data <=  16;
			when 280 => sin_inv_data <=  16;
			when 281 => sin_inv_data <=  16;
			when 282 => sin_inv_data <=  16;
			when 283 => sin_inv_data <=  16;
			when 284 => sin_inv_data <=  16;
			when 285 => sin_inv_data <=  17;
			when 286 => sin_inv_data <=  17;
			when 287 => sin_inv_data <=  17;
			when 288 => sin_inv_data <=  17;
			when 289 => sin_inv_data <=  17;
			when 290 => sin_inv_data <=  17;
			when 291 => sin_inv_data <=  17;
			when 292 => sin_inv_data <=  17;
			when 293 => sin_inv_data <=  17;
			when 294 => sin_inv_data <=  17;
			when 295 => sin_inv_data <=  17;
			when 296 => sin_inv_data <=  17;
			when 297 => sin_inv_data <=  17;
			when 298 => sin_inv_data <=  17;
			when 299 => sin_inv_data <=  17;
			when 300 => sin_inv_data <=  17;
			when 301 => sin_inv_data <=  18;
			when 302 => sin_inv_data <=  18;
			when 303 => sin_inv_data <=  18;
			when 304 => sin_inv_data <=  18;
			when 305 => sin_inv_data <=  18;
			when 306 => sin_inv_data <=  18;
			when 307 => sin_inv_data <=  18;
			when 308 => sin_inv_data <=  18;
			when 309 => sin_inv_data <=  18;
			when 310 => sin_inv_data <=  18;
			when 311 => sin_inv_data <=  18;
			when 312 => sin_inv_data <=  18;
			when 313 => sin_inv_data <=  18;
			when 314 => sin_inv_data <=  18;
			when 315 => sin_inv_data <=  18;
			when 316 => sin_inv_data <=  18;
			when 317 => sin_inv_data <=  18;
			when 318 => sin_inv_data <=  19;
			when 319 => sin_inv_data <=  19;
			when 320 => sin_inv_data <=  19;
			when 321 => sin_inv_data <=  19;
			when 322 => sin_inv_data <=  19;
			when 323 => sin_inv_data <=  19;
			when 324 => sin_inv_data <=  19;
			when 325 => sin_inv_data <=  19;
			when 326 => sin_inv_data <=  19;
			when 327 => sin_inv_data <=  19;
			when 328 => sin_inv_data <=  19;
			when 329 => sin_inv_data <=  19;
			when 330 => sin_inv_data <=  19;
			when 331 => sin_inv_data <=  19;
			when 332 => sin_inv_data <=  19;
			when 333 => sin_inv_data <=  19;
			when 334 => sin_inv_data <=  20;
			when 335 => sin_inv_data <=  20;
			when 336 => sin_inv_data <=  20;
			when 337 => sin_inv_data <=  20;
			when 338 => sin_inv_data <=  20;
			when 339 => sin_inv_data <=  20;
			when 340 => sin_inv_data <=  20;
			when 341 => sin_inv_data <=  20;
			when 342 => sin_inv_data <=  20;
			when 343 => sin_inv_data <=  20;
			when 344 => sin_inv_data <=  20;
			when 345 => sin_inv_data <=  20;
			when 346 => sin_inv_data <=  20;
			when 347 => sin_inv_data <=  20;
			when 348 => sin_inv_data <=  20;
			when 349 => sin_inv_data <=  20;
			when 350 => sin_inv_data <=  20;
			when 351 => sin_inv_data <=  21;
			when 352 => sin_inv_data <=  21;
			when 353 => sin_inv_data <=  21;
			when 354 => sin_inv_data <=  21;
			when 355 => sin_inv_data <=  21;
			when 356 => sin_inv_data <=  21;
			when 357 => sin_inv_data <=  21;
			when 358 => sin_inv_data <=  21;
			when 359 => sin_inv_data <=  21;
			when 360 => sin_inv_data <=  21;
			when 361 => sin_inv_data <=  21;
			when 362 => sin_inv_data <=  21;
			when 363 => sin_inv_data <=  21;
			when 364 => sin_inv_data <=  21;
			when 365 => sin_inv_data <=  21;
			when 366 => sin_inv_data <=  21;
			when 367 => sin_inv_data <=  22;
			when 368 => sin_inv_data <=  22;
			when 369 => sin_inv_data <=  22;
			when 370 => sin_inv_data <=  22;
			when 371 => sin_inv_data <=  22;
			when 372 => sin_inv_data <=  22;
			when 373 => sin_inv_data <=  22;
			when 374 => sin_inv_data <=  22;
			when 375 => sin_inv_data <=  22;
			when 376 => sin_inv_data <=  22;
			when 377 => sin_inv_data <=  22;
			when 378 => sin_inv_data <=  22;
			when 379 => sin_inv_data <=  22;
			when 380 => sin_inv_data <=  22;
			when 381 => sin_inv_data <=  22;
			when 382 => sin_inv_data <=  22;
			when 383 => sin_inv_data <=  23;
			when 384 => sin_inv_data <=  23;
			when 385 => sin_inv_data <=  23;
			when 386 => sin_inv_data <=  23;
			when 387 => sin_inv_data <=  23;
			when 388 => sin_inv_data <=  23;
			when 389 => sin_inv_data <=  23;
			when 390 => sin_inv_data <=  23;
			when 391 => sin_inv_data <=  23;
			when 392 => sin_inv_data <=  23;
			when 393 => sin_inv_data <=  23;
			when 394 => sin_inv_data <=  23;
			when 395 => sin_inv_data <=  23;
			when 396 => sin_inv_data <=  23;
			when 397 => sin_inv_data <=  23;
			when 398 => sin_inv_data <=  23;
			when 399 => sin_inv_data <=  24;
			when 400 => sin_inv_data <=  24;
			when 401 => sin_inv_data <=  24;
			when 402 => sin_inv_data <=  24;
			when 403 => sin_inv_data <=  24;
			when 404 => sin_inv_data <=  24;
			when 405 => sin_inv_data <=  24;
			when 406 => sin_inv_data <=  24;
			when 407 => sin_inv_data <=  24;
			when 408 => sin_inv_data <=  24;
			when 409 => sin_inv_data <=  24;
			when 410 => sin_inv_data <=  24;
			when 411 => sin_inv_data <=  24;
			when 412 => sin_inv_data <=  24;
			when 413 => sin_inv_data <=  24;
			when 414 => sin_inv_data <=  24;
			when 415 => sin_inv_data <=  25;
			when 416 => sin_inv_data <=  25;
			when 417 => sin_inv_data <=  25;
			when 418 => sin_inv_data <=  25;
			when 419 => sin_inv_data <=  25;
			when 420 => sin_inv_data <=  25;
			when 421 => sin_inv_data <=  25;
			when 422 => sin_inv_data <=  25;
			when 423 => sin_inv_data <=  25;
			when 424 => sin_inv_data <=  25;
			when 425 => sin_inv_data <=  25;
			when 426 => sin_inv_data <=  25;
			when 427 => sin_inv_data <=  25;
			when 428 => sin_inv_data <=  25;
			when 429 => sin_inv_data <=  25;
			when 430 => sin_inv_data <=  25;
			when 431 => sin_inv_data <=  26;
			when 432 => sin_inv_data <=  26;
			when 433 => sin_inv_data <=  26;
			when 434 => sin_inv_data <=  26;
			when 435 => sin_inv_data <=  26;
			when 436 => sin_inv_data <=  26;
			when 437 => sin_inv_data <=  26;
			when 438 => sin_inv_data <=  26;
			when 439 => sin_inv_data <=  26;
			when 440 => sin_inv_data <=  26;
			when 441 => sin_inv_data <=  26;
			when 442 => sin_inv_data <=  26;
			when 443 => sin_inv_data <=  26;
			when 444 => sin_inv_data <=  26;
			when 445 => sin_inv_data <=  26;
			when 446 => sin_inv_data <=  26;
			when 447 => sin_inv_data <=  27;
			when 448 => sin_inv_data <=  27;
			when 449 => sin_inv_data <=  27;
			when 450 => sin_inv_data <=  27;
			when 451 => sin_inv_data <=  27;
			when 452 => sin_inv_data <=  27;
			when 453 => sin_inv_data <=  27;
			when 454 => sin_inv_data <=  27;
			when 455 => sin_inv_data <=  27;
			when 456 => sin_inv_data <=  27;
			when 457 => sin_inv_data <=  27;
			when 458 => sin_inv_data <=  27;
			when 459 => sin_inv_data <=  27;
			when 460 => sin_inv_data <=  27;
			when 461 => sin_inv_data <=  27;
			when 462 => sin_inv_data <=  28;
			when 463 => sin_inv_data <=  28;
			when 464 => sin_inv_data <=  28;
			when 465 => sin_inv_data <=  28;
			when 466 => sin_inv_data <=  28;
			when 467 => sin_inv_data <=  28;
			when 468 => sin_inv_data <=  28;
			when 469 => sin_inv_data <=  28;
			when 470 => sin_inv_data <=  28;
			when 471 => sin_inv_data <=  28;
			when 472 => sin_inv_data <=  28;
			when 473 => sin_inv_data <=  28;
			when 474 => sin_inv_data <=  28;
			when 475 => sin_inv_data <=  28;
			when 476 => sin_inv_data <=  28;
			when 477 => sin_inv_data <=  28;
			when 478 => sin_inv_data <=  29;
			when 479 => sin_inv_data <=  29;
			when 480 => sin_inv_data <=  29;
			when 481 => sin_inv_data <=  29;
			when 482 => sin_inv_data <=  29;
			when 483 => sin_inv_data <=  29;
			when 484 => sin_inv_data <=  29;
			when 485 => sin_inv_data <=  29;
			when 486 => sin_inv_data <=  29;
			when 487 => sin_inv_data <=  29;
			when 488 => sin_inv_data <=  29;
			when 489 => sin_inv_data <=  29;
			when 490 => sin_inv_data <=  29;
			when 491 => sin_inv_data <=  29;
			when 492 => sin_inv_data <=  29;
			when 493 => sin_inv_data <=  30;
			when 494 => sin_inv_data <=  30;
			when 495 => sin_inv_data <=  30;
			when 496 => sin_inv_data <=  30;
			when 497 => sin_inv_data <=  30;
			when 498 => sin_inv_data <=  30;
			when 499 => sin_inv_data <=  30;
			when 500 => sin_inv_data <=  30;
			when 501 => sin_inv_data <=  30;
			when 502 => sin_inv_data <=  30;
			when 503 => sin_inv_data <=  30;
			when 504 => sin_inv_data <=  30;
			when 505 => sin_inv_data <=  30;
			when 506 => sin_inv_data <=  30;
			when 507 => sin_inv_data <=  30;
			when 508 => sin_inv_data <=  31;
			when 509 => sin_inv_data <=  31;
			when 510 => sin_inv_data <=  31;
			when 511 => sin_inv_data <=  31;
			when 512 => sin_inv_data <=  31;
			when 513 => sin_inv_data <=  31;
			when 514 => sin_inv_data <=  31;
			when 515 => sin_inv_data <=  31;
			when 516 => sin_inv_data <=  31;
			when 517 => sin_inv_data <=  31;
			when 518 => sin_inv_data <=  31;
			when 519 => sin_inv_data <=  31;
			when 520 => sin_inv_data <=  31;
			when 521 => sin_inv_data <=  31;
			when 522 => sin_inv_data <=  31;
			when 523 => sin_inv_data <=  32;
			when 524 => sin_inv_data <=  32;
			when 525 => sin_inv_data <=  32;
			when 526 => sin_inv_data <=  32;
			when 527 => sin_inv_data <=  32;
			when 528 => sin_inv_data <=  32;
			when 529 => sin_inv_data <=  32;
			when 530 => sin_inv_data <=  32;
			when 531 => sin_inv_data <=  32;
			when 532 => sin_inv_data <=  32;
			when 533 => sin_inv_data <=  32;
			when 534 => sin_inv_data <=  32;
			when 535 => sin_inv_data <=  32;
			when 536 => sin_inv_data <=  32;
			when 537 => sin_inv_data <=  32;
			when 538 => sin_inv_data <=  33;
			when 539 => sin_inv_data <=  33;
			when 540 => sin_inv_data <=  33;
			when 541 => sin_inv_data <=  33;
			when 542 => sin_inv_data <=  33;
			when 543 => sin_inv_data <=  33;
			when 544 => sin_inv_data <=  33;
			when 545 => sin_inv_data <=  33;
			when 546 => sin_inv_data <=  33;
			when 547 => sin_inv_data <=  33;
			when 548 => sin_inv_data <=  33;
			when 549 => sin_inv_data <=  33;
			when 550 => sin_inv_data <=  33;
			when 551 => sin_inv_data <=  33;
			when 552 => sin_inv_data <=  34;
			when 553 => sin_inv_data <=  34;
			when 554 => sin_inv_data <=  34;
			when 555 => sin_inv_data <=  34;
			when 556 => sin_inv_data <=  34;
			when 557 => sin_inv_data <=  34;
			when 558 => sin_inv_data <=  34;
			when 559 => sin_inv_data <=  34;
			when 560 => sin_inv_data <=  34;
			when 561 => sin_inv_data <=  34;
			when 562 => sin_inv_data <=  34;
			when 563 => sin_inv_data <=  34;
			when 564 => sin_inv_data <=  34;
			when 565 => sin_inv_data <=  34;
			when 566 => sin_inv_data <=  34;
			when 567 => sin_inv_data <=  35;
			when 568 => sin_inv_data <=  35;
			when 569 => sin_inv_data <=  35;
			when 570 => sin_inv_data <=  35;
			when 571 => sin_inv_data <=  35;
			when 572 => sin_inv_data <=  35;
			when 573 => sin_inv_data <=  35;
			when 574 => sin_inv_data <=  35;
			when 575 => sin_inv_data <=  35;
			when 576 => sin_inv_data <=  35;
			when 577 => sin_inv_data <=  35;
			when 578 => sin_inv_data <=  35;
			when 579 => sin_inv_data <=  35;
			when 580 => sin_inv_data <=  35;
			when 581 => sin_inv_data <=  36;
			when 582 => sin_inv_data <=  36;
			when 583 => sin_inv_data <=  36;
			when 584 => sin_inv_data <=  36;
			when 585 => sin_inv_data <=  36;
			when 586 => sin_inv_data <=  36;
			when 587 => sin_inv_data <=  36;
			when 588 => sin_inv_data <=  36;
			when 589 => sin_inv_data <=  36;
			when 590 => sin_inv_data <=  36;
			when 591 => sin_inv_data <=  36;
			when 592 => sin_inv_data <=  36;
			when 593 => sin_inv_data <=  36;
			when 594 => sin_inv_data <=  36;
			when 595 => sin_inv_data <=  37;
			when 596 => sin_inv_data <=  37;
			when 597 => sin_inv_data <=  37;
			when 598 => sin_inv_data <=  37;
			when 599 => sin_inv_data <=  37;
			when 600 => sin_inv_data <=  37;
			when 601 => sin_inv_data <=  37;
			when 602 => sin_inv_data <=  37;
			when 603 => sin_inv_data <=  37;
			when 604 => sin_inv_data <=  37;
			when 605 => sin_inv_data <=  37;
			when 606 => sin_inv_data <=  37;
			when 607 => sin_inv_data <=  37;
			when 608 => sin_inv_data <=  37;
			when 609 => sin_inv_data <=  38;
			when 610 => sin_inv_data <=  38;
			when 611 => sin_inv_data <=  38;
			when 612 => sin_inv_data <=  38;
			when 613 => sin_inv_data <=  38;
			when 614 => sin_inv_data <=  38;
			when 615 => sin_inv_data <=  38;
			when 616 => sin_inv_data <=  38;
			when 617 => sin_inv_data <=  38;
			when 618 => sin_inv_data <=  38;
			when 619 => sin_inv_data <=  38;
			when 620 => sin_inv_data <=  38;
			when 621 => sin_inv_data <=  38;
			when 622 => sin_inv_data <=  38;
			when 623 => sin_inv_data <=  39;
			when 624 => sin_inv_data <=  39;
			when 625 => sin_inv_data <=  39;
			when 626 => sin_inv_data <=  39;
			when 627 => sin_inv_data <=  39;
			when 628 => sin_inv_data <=  39;
			when 629 => sin_inv_data <=  39;
			when 630 => sin_inv_data <=  39;
			when 631 => sin_inv_data <=  39;
			when 632 => sin_inv_data <=  39;
			when 633 => sin_inv_data <=  39;
			when 634 => sin_inv_data <=  39;
			when 635 => sin_inv_data <=  39;
			when 636 => sin_inv_data <=  39;
			when 637 => sin_inv_data <=  40;
			when 638 => sin_inv_data <=  40;
			when 639 => sin_inv_data <=  40;
			when 640 => sin_inv_data <=  40;
			when 641 => sin_inv_data <=  40;
			when 642 => sin_inv_data <=  40;
			when 643 => sin_inv_data <=  40;
			when 644 => sin_inv_data <=  40;
			when 645 => sin_inv_data <=  40;
			when 646 => sin_inv_data <=  40;
			when 647 => sin_inv_data <=  40;
			when 648 => sin_inv_data <=  40;
			when 649 => sin_inv_data <=  40;
			when 650 => sin_inv_data <=  41;
			when 651 => sin_inv_data <=  41;
			when 652 => sin_inv_data <=  41;
			when 653 => sin_inv_data <=  41;
			when 654 => sin_inv_data <=  41;
			when 655 => sin_inv_data <=  41;
			when 656 => sin_inv_data <=  41;
			when 657 => sin_inv_data <=  41;
			when 658 => sin_inv_data <=  41;
			when 659 => sin_inv_data <=  41;
			when 660 => sin_inv_data <=  41;
			when 661 => sin_inv_data <=  41;
			when 662 => sin_inv_data <=  41;
			when 663 => sin_inv_data <=  42;
			when 664 => sin_inv_data <=  42;
			when 665 => sin_inv_data <=  42;
			when 666 => sin_inv_data <=  42;
			when 667 => sin_inv_data <=  42;
			when 668 => sin_inv_data <=  42;
			when 669 => sin_inv_data <=  42;
			when 670 => sin_inv_data <=  42;
			when 671 => sin_inv_data <=  42;
			when 672 => sin_inv_data <=  42;
			when 673 => sin_inv_data <=  42;
			when 674 => sin_inv_data <=  42;
			when 675 => sin_inv_data <=  42;
			when 676 => sin_inv_data <=  43;
			when 677 => sin_inv_data <=  43;
			when 678 => sin_inv_data <=  43;
			when 679 => sin_inv_data <=  43;
			when 680 => sin_inv_data <=  43;
			when 681 => sin_inv_data <=  43;
			when 682 => sin_inv_data <=  43;
			when 683 => sin_inv_data <=  43;
			when 684 => sin_inv_data <=  43;
			when 685 => sin_inv_data <=  43;
			when 686 => sin_inv_data <=  43;
			when 687 => sin_inv_data <=  43;
			when 688 => sin_inv_data <=  43;
			when 689 => sin_inv_data <=  44;
			when 690 => sin_inv_data <=  44;
			when 691 => sin_inv_data <=  44;
			when 692 => sin_inv_data <=  44;
			when 693 => sin_inv_data <=  44;
			when 694 => sin_inv_data <=  44;
			when 695 => sin_inv_data <=  44;
			when 696 => sin_inv_data <=  44;
			when 697 => sin_inv_data <=  44;
			when 698 => sin_inv_data <=  44;
			when 699 => sin_inv_data <=  44;
			when 700 => sin_inv_data <=  44;
			when 701 => sin_inv_data <=  45;
			when 702 => sin_inv_data <=  45;
			when 703 => sin_inv_data <=  45;
			when 704 => sin_inv_data <=  45;
			when 705 => sin_inv_data <=  45;
			when 706 => sin_inv_data <=  45;
			when 707 => sin_inv_data <=  45;
			when 708 => sin_inv_data <=  45;
			when 709 => sin_inv_data <=  45;
			when 710 => sin_inv_data <=  45;
			when 711 => sin_inv_data <=  45;
			when 712 => sin_inv_data <=  45;
			when 713 => sin_inv_data <=  45;
			when 714 => sin_inv_data <=  46;
			when 715 => sin_inv_data <=  46;
			when 716 => sin_inv_data <=  46;
			when 717 => sin_inv_data <=  46;
			when 718 => sin_inv_data <=  46;
			when 719 => sin_inv_data <=  46;
			when 720 => sin_inv_data <=  46;
			when 721 => sin_inv_data <=  46;
			when 722 => sin_inv_data <=  46;
			when 723 => sin_inv_data <=  46;
			when 724 => sin_inv_data <=  46;
			when 725 => sin_inv_data <=  46;
			when 726 => sin_inv_data <=  47;
			when 727 => sin_inv_data <=  47;
			when 728 => sin_inv_data <=  47;
			when 729 => sin_inv_data <=  47;
			when 730 => sin_inv_data <=  47;
			when 731 => sin_inv_data <=  47;
			when 732 => sin_inv_data <=  47;
			when 733 => sin_inv_data <=  47;
			when 734 => sin_inv_data <=  47;
			when 735 => sin_inv_data <=  47;
			when 736 => sin_inv_data <=  47;
			when 737 => sin_inv_data <=  47;
			when 738 => sin_inv_data <=  48;
			when 739 => sin_inv_data <=  48;
			when 740 => sin_inv_data <=  48;
			when 741 => sin_inv_data <=  48;
			when 742 => sin_inv_data <=  48;
			when 743 => sin_inv_data <=  48;
			when 744 => sin_inv_data <=  48;
			when 745 => sin_inv_data <=  48;
			when 746 => sin_inv_data <=  48;
			when 747 => sin_inv_data <=  48;
			when 748 => sin_inv_data <=  48;
			when 749 => sin_inv_data <=  49;
			when 750 => sin_inv_data <=  49;
			when 751 => sin_inv_data <=  49;
			when 752 => sin_inv_data <=  49;
			when 753 => sin_inv_data <=  49;
			when 754 => sin_inv_data <=  49;
			when 755 => sin_inv_data <=  49;
			when 756 => sin_inv_data <=  49;
			when 757 => sin_inv_data <=  49;
			when 758 => sin_inv_data <=  49;
			when 759 => sin_inv_data <=  49;
			when 760 => sin_inv_data <=  49;
			when 761 => sin_inv_data <=  50;
			when 762 => sin_inv_data <=  50;
			when 763 => sin_inv_data <=  50;
			when 764 => sin_inv_data <=  50;
			when 765 => sin_inv_data <=  50;
			when 766 => sin_inv_data <=  50;
			when 767 => sin_inv_data <=  50;
			when 768 => sin_inv_data <=  50;
			when 769 => sin_inv_data <=  50;
			when 770 => sin_inv_data <=  50;
			when 771 => sin_inv_data <=  50;
			when 772 => sin_inv_data <=  51;
			when 773 => sin_inv_data <=  51;
			when 774 => sin_inv_data <=  51;
			when 775 => sin_inv_data <=  51;
			when 776 => sin_inv_data <=  51;
			when 777 => sin_inv_data <=  51;
			when 778 => sin_inv_data <=  51;
			when 779 => sin_inv_data <=  51;
			when 780 => sin_inv_data <=  51;
			when 781 => sin_inv_data <=  51;
			when 782 => sin_inv_data <=  51;
			when 783 => sin_inv_data <=  52;
			when 784 => sin_inv_data <=  52;
			when 785 => sin_inv_data <=  52;
			when 786 => sin_inv_data <=  52;
			when 787 => sin_inv_data <=  52;
			when 788 => sin_inv_data <=  52;
			when 789 => sin_inv_data <=  52;
			when 790 => sin_inv_data <=  52;
			when 791 => sin_inv_data <=  52;
			when 792 => sin_inv_data <=  52;
			when 793 => sin_inv_data <=  52;
			when 794 => sin_inv_data <=  53;
			when 795 => sin_inv_data <=  53;
			when 796 => sin_inv_data <=  53;
			when 797 => sin_inv_data <=  53;
			when 798 => sin_inv_data <=  53;
			when 799 => sin_inv_data <=  53;
			when 800 => sin_inv_data <=  53;
			when 801 => sin_inv_data <=  53;
			when 802 => sin_inv_data <=  53;
			when 803 => sin_inv_data <=  53;
			when 804 => sin_inv_data <=  54;
			when 805 => sin_inv_data <=  54;
			when 806 => sin_inv_data <=  54;
			when 807 => sin_inv_data <=  54;
			when 808 => sin_inv_data <=  54;
			when 809 => sin_inv_data <=  54;
			when 810 => sin_inv_data <=  54;
			when 811 => sin_inv_data <=  54;
			when 812 => sin_inv_data <=  54;
			when 813 => sin_inv_data <=  54;
			when 814 => sin_inv_data <=  54;
			when 815 => sin_inv_data <=  55;
			when 816 => sin_inv_data <=  55;
			when 817 => sin_inv_data <=  55;
			when 818 => sin_inv_data <=  55;
			when 819 => sin_inv_data <=  55;
			when 820 => sin_inv_data <=  55;
			when 821 => sin_inv_data <=  55;
			when 822 => sin_inv_data <=  55;
			when 823 => sin_inv_data <=  55;
			when 824 => sin_inv_data <=  55;
			when 825 => sin_inv_data <=  56;
			when 826 => sin_inv_data <=  56;
			when 827 => sin_inv_data <=  56;
			when 828 => sin_inv_data <=  56;
			when 829 => sin_inv_data <=  56;
			when 830 => sin_inv_data <=  56;
			when 831 => sin_inv_data <=  56;
			when 832 => sin_inv_data <=  56;
			when 833 => sin_inv_data <=  56;
			when 834 => sin_inv_data <=  57;
			when 835 => sin_inv_data <=  57;
			when 836 => sin_inv_data <=  57;
			when 837 => sin_inv_data <=  57;
			when 838 => sin_inv_data <=  57;
			when 839 => sin_inv_data <=  57;
			when 840 => sin_inv_data <=  57;
			when 841 => sin_inv_data <=  57;
			when 842 => sin_inv_data <=  57;
			when 843 => sin_inv_data <=  57;
			when 844 => sin_inv_data <=  58;
			when 845 => sin_inv_data <=  58;
			when 846 => sin_inv_data <=  58;
			when 847 => sin_inv_data <=  58;
			when 848 => sin_inv_data <=  58;
			when 849 => sin_inv_data <=  58;
			when 850 => sin_inv_data <=  58;
			when 851 => sin_inv_data <=  58;
			when 852 => sin_inv_data <=  58;
			when 853 => sin_inv_data <=  59;
			when 854 => sin_inv_data <=  59;
			when 855 => sin_inv_data <=  59;
			when 856 => sin_inv_data <=  59;
			when 857 => sin_inv_data <=  59;
			when 858 => sin_inv_data <=  59;
			when 859 => sin_inv_data <=  59;
			when 860 => sin_inv_data <=  59;
			when 861 => sin_inv_data <=  59;
			when 862 => sin_inv_data <=  60;
			when 863 => sin_inv_data <=  60;
			when 864 => sin_inv_data <=  60;
			when 865 => sin_inv_data <=  60;
			when 866 => sin_inv_data <=  60;
			when 867 => sin_inv_data <=  60;
			when 868 => sin_inv_data <=  60;
			when 869 => sin_inv_data <=  60;
			when 870 => sin_inv_data <=  60;
			when 871 => sin_inv_data <=  61;
			when 872 => sin_inv_data <=  61;
			when 873 => sin_inv_data <=  61;
			when 874 => sin_inv_data <=  61;
			when 875 => sin_inv_data <=  61;
			when 876 => sin_inv_data <=  61;
			when 877 => sin_inv_data <=  61;
			when 878 => sin_inv_data <=  61;
			when 879 => sin_inv_data <=  62;
			when 880 => sin_inv_data <=  62;
			when 881 => sin_inv_data <=  62;
			when 882 => sin_inv_data <=  62;
			when 883 => sin_inv_data <=  62;
			when 884 => sin_inv_data <=  62;
			when 885 => sin_inv_data <=  62;
			when 886 => sin_inv_data <=  62;
			when 887 => sin_inv_data <=  62;
			when 888 => sin_inv_data <=  63;
			when 889 => sin_inv_data <=  63;
			when 890 => sin_inv_data <=  63;
			when 891 => sin_inv_data <=  63;
			when 892 => sin_inv_data <=  63;
			when 893 => sin_inv_data <=  63;
			when 894 => sin_inv_data <=  63;
			when 895 => sin_inv_data <=  64;
			when 896 => sin_inv_data <=  64;
			when 897 => sin_inv_data <=  64;
			when 898 => sin_inv_data <=  64;
			when 899 => sin_inv_data <=  64;
			when 900 => sin_inv_data <=  64;
			when 901 => sin_inv_data <=  64;
			when 902 => sin_inv_data <=  64;
			when 903 => sin_inv_data <=  65;
			when 904 => sin_inv_data <=  65;
			when 905 => sin_inv_data <=  65;
			when 906 => sin_inv_data <=  65;
			when 907 => sin_inv_data <=  65;
			when 908 => sin_inv_data <=  65;
			when 909 => sin_inv_data <=  65;
			when 910 => sin_inv_data <=  66;
			when 911 => sin_inv_data <=  66;
			when 912 => sin_inv_data <=  66;
			when 913 => sin_inv_data <=  66;
			when 914 => sin_inv_data <=  66;
			when 915 => sin_inv_data <=  66;
			when 916 => sin_inv_data <=  66;
			when 917 => sin_inv_data <=  66;
			when 918 => sin_inv_data <=  67;
			when 919 => sin_inv_data <=  67;
			when 920 => sin_inv_data <=  67;
			when 921 => sin_inv_data <=  67;
			when 922 => sin_inv_data <=  67;
			when 923 => sin_inv_data <=  67;
			when 924 => sin_inv_data <=  68;
			when 925 => sin_inv_data <=  68;
			when 926 => sin_inv_data <=  68;
			when 927 => sin_inv_data <=  68;
			when 928 => sin_inv_data <=  68;
			when 929 => sin_inv_data <=  68;
			when 930 => sin_inv_data <=  68;
			when 931 => sin_inv_data <=  69;
			when 932 => sin_inv_data <=  69;
			when 933 => sin_inv_data <=  69;
			when 934 => sin_inv_data <=  69;
			when 935 => sin_inv_data <=  69;
			when 936 => sin_inv_data <=  69;
			when 937 => sin_inv_data <=  70;
			when 938 => sin_inv_data <=  70;
			when 939 => sin_inv_data <=  70;
			when 940 => sin_inv_data <=  70;
			when 941 => sin_inv_data <=  70;
			when 942 => sin_inv_data <=  70;
			when 943 => sin_inv_data <=  71;
			when 944 => sin_inv_data <=  71;
			when 945 => sin_inv_data <=  71;
			when 946 => sin_inv_data <=  71;
			when 947 => sin_inv_data <=  71;
			when 948 => sin_inv_data <=  71;
			when 949 => sin_inv_data <=  72;
			when 950 => sin_inv_data <=  72;
			when 951 => sin_inv_data <=  72;
			when 952 => sin_inv_data <=  72;
			when 953 => sin_inv_data <=  72;
			when 954 => sin_inv_data <=  73;
			when 955 => sin_inv_data <=  73;
			when 956 => sin_inv_data <=  73;
			when 957 => sin_inv_data <=  73;
			when 958 => sin_inv_data <=  73;
			when 959 => sin_inv_data <=  74;
			when 960 => sin_inv_data <=  74;
			when 961 => sin_inv_data <=  74;
			when 962 => sin_inv_data <=  74;
			when 963 => sin_inv_data <=  74;
			when 964 => sin_inv_data <=  75;
			when 965 => sin_inv_data <=  75;
			when 966 => sin_inv_data <=  75;
			when 967 => sin_inv_data <=  75;
			when 968 => sin_inv_data <=  75;
			when 969 => sin_inv_data <=  76;
			when 970 => sin_inv_data <=  76;
			when 971 => sin_inv_data <=  76;
			when 972 => sin_inv_data <=  76;
			when 973 => sin_inv_data <=  77;
			when 974 => sin_inv_data <=  77;
			when 975 => sin_inv_data <=  77;
			when 976 => sin_inv_data <=  77;
			when 977 => sin_inv_data <=  78;
			when 978 => sin_inv_data <=  78;
			when 979 => sin_inv_data <=  78;
			when 980 => sin_inv_data <=  79;
			when 981 => sin_inv_data <=  79;
			when 982 => sin_inv_data <=  79;
			when 983 => sin_inv_data <=  79;
			when 984 => sin_inv_data <=  80;
			when 985 => sin_inv_data <=  80;
			when 986 => sin_inv_data <=  80;
			when 987 => sin_inv_data <=  81;
			when 988 => sin_inv_data <=  81;
			when 989 => sin_inv_data <=  81;
			when 990 => sin_inv_data <=  82;
			when 991 => sin_inv_data <=  82;
			when 992 => sin_inv_data <=  83;
			when 993 => sin_inv_data <=  83;
			when 994 => sin_inv_data <=  84;
			when 995 => sin_inv_data <=  84;
			when 996 => sin_inv_data <=  85;
			when 997 => sin_inv_data <=  86;
			when 998 => sin_inv_data <=  86;
			when 999 => sin_inv_data <=  87;
			when 1000 => sin_inv_data <=  90;

      when others       => null;
      end case;
	
		
		end if;
   end if;
end process;


end rtl;
