
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sincos_lut is
port
(
   clk               :  IN  std_logic;
	reset 				: 	IN STD_LOGIC;
	clk_50				: 	IN STD_LOGIC;
	avs_s0_address		: 	IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	avs_s0_read			: 	IN STD_LOGIC;
	avs_s0_write		: 	IN STD_LOGIC;
	avs_s0_readdata	: 	OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
	avs_s0_writedata	: 	IN STD_LOGIC_VECTOR(31 DOWNTO 0)

);

end sincos_lut;


architecture rtl of sincos_lut is
   signal theta           : std_logic_vector(31 downto 0); --11 downto 0
   signal sin_data        : signed(31 downto 0);
   signal cos_data        : signed(31 downto 0);
   --signal theta_int     : integer range 0 to 4095 := 0;
   signal sin_data_int    : signed(31 downto 0);
   signal cos_data_int    : signed(31 downto 0);
   signal reset_n         : std_logic;
   signal clk_en          : std_logic;signal led : std_logic_vector(7 downto 0); 

begin



   AV_READ: PROCESS(clk)
	BEGIN
		IF rising_edge(clk) THEN
			IF (reset='1') THEN
				avs_s0_readdata <= x"00000000";
				ELSIF (avs_s0_read='1') THEN
					IF (avs_s0_address = x"00" )THEN
						avs_s0_readdata 	<=		std_logic_vector(sin_data(31 downto 0)) AND x"FFFFFFFF"; 
					 ELSIF (avs_s0_address = x"01") THEN
						avs_s0_readdata 	<=		std_logic_vector(cos_data(31 downto 0)) AND x"FFFFFFFF"; 
					
					ELSE avs_s0_readdata <= x"0000ffff";
				END IF;		
			END IF;
		END IF;
	END PROCESS;
		 
	  AV_WRITE: PROCESS(clk)
	  --variable read_data : std_logic_vector(31 downto 0):= x"00000000";

	  BEGIN
        IF rising_edge(clk) THEN
            IF (reset='1') THEN
                led <= "00001111";
            ELSIF (avs_s0_write='1') THEN               
					 IF (avs_s0_address = x"00" )THEN
                    theta 				<= avs_s0_writedata(31 downto 0); --start
 					 ELSIF (avs_s0_address = x"01") THEN
                    clk_en 		   <= avs_s0_writedata(0); --pressure
						  reset_n         <= NOT(clk_en);
					 ELSE led 						<= "11110000";
					 END IF; 
            END IF;
        END IF;
	  END PROCESS;	


sin_cos_lut: process(clk_50)
	variable theta_int  : integer range 0 to 4095 := 0;
	begin
   if(reset_n = '1')then
       sin_data_int <= to_signed(3500,32); 
       cos_data_int <= to_signed(3500,32);
   elsif(rising_edge(clk_50)) then
      if clk_en = '1' then
         theta_int := to_integer(unsigned(theta));

         sin_data <= sin_data_int;
         cos_data <= cos_data_int;

         case theta_int is
				when 0 => sin_data_int <= to_signed(0,32); cos_data_int <= to_signed(1000,32);
				when 1 => sin_data_int <= to_signed(2,32); cos_data_int <= to_signed(1000,32);
				when 2 => sin_data_int <= to_signed(3,32); cos_data_int <= to_signed(1000,32);
				when 3 => sin_data_int <= to_signed(5,32); cos_data_int <= to_signed(1000,32);
				when 4 => sin_data_int <= to_signed(6,32); cos_data_int <= to_signed(1000,32);
				when 5 => sin_data_int <= to_signed(8,32); cos_data_int <= to_signed(1000,32);
				when 6 => sin_data_int <= to_signed(9,32); cos_data_int <= to_signed(1000,32);
				when 7 => sin_data_int <= to_signed(11,32); cos_data_int <= to_signed(1000,32);
				when 8 => sin_data_int <= to_signed(12,32); cos_data_int <= to_signed(1000,32);
				when 9 => sin_data_int <= to_signed(14,32); cos_data_int <= to_signed(1000,32);
				when 10 => sin_data_int <= to_signed(15,32); cos_data_int <= to_signed(1000,32);
				when 11 => sin_data_int <= to_signed(17,32); cos_data_int <= to_signed(1000,32);
				when 12 => sin_data_int <= to_signed(18,32); cos_data_int <= to_signed(1000,32);
				when 13 => sin_data_int <= to_signed(20,32); cos_data_int <= to_signed(1000,32);
				when 14 => sin_data_int <= to_signed(21,32); cos_data_int <= to_signed(1000,32);
				when 15 => sin_data_int <= to_signed(23,32); cos_data_int <= to_signed(1000,32);
				when 16 => sin_data_int <= to_signed(25,32); cos_data_int <= to_signed(1000,32);
				when 17 => sin_data_int <= to_signed(26,32); cos_data_int <= to_signed(1000,32);
				when 18 => sin_data_int <= to_signed(28,32); cos_data_int <= to_signed(1000,32);
				when 19 => sin_data_int <= to_signed(29,32); cos_data_int <= to_signed(1000,32);
				when 20 => sin_data_int <= to_signed(31,32); cos_data_int <= to_signed(999,32);
				when 21 => sin_data_int <= to_signed(32,32); cos_data_int <= to_signed(999,32);
				when 22 => sin_data_int <= to_signed(34,32); cos_data_int <= to_signed(999,32);
				when 23 => sin_data_int <= to_signed(35,32); cos_data_int <= to_signed(999,32);
				when 24 => sin_data_int <= to_signed(37,32); cos_data_int <= to_signed(999,32);
				when 25 => sin_data_int <= to_signed(38,32); cos_data_int <= to_signed(999,32);
				when 26 => sin_data_int <= to_signed(40,32); cos_data_int <= to_signed(999,32);
				when 27 => sin_data_int <= to_signed(41,32); cos_data_int <= to_signed(999,32);
				when 28 => sin_data_int <= to_signed(43,32); cos_data_int <= to_signed(999,32);
				when 29 => sin_data_int <= to_signed(44,32); cos_data_int <= to_signed(999,32);
				when 30 => sin_data_int <= to_signed(46,32); cos_data_int <= to_signed(999,32);
				when 31 => sin_data_int <= to_signed(48,32); cos_data_int <= to_signed(999,32);
				when 32 => sin_data_int <= to_signed(49,32); cos_data_int <= to_signed(999,32);
				when 33 => sin_data_int <= to_signed(51,32); cos_data_int <= to_signed(999,32);
				when 34 => sin_data_int <= to_signed(52,32); cos_data_int <= to_signed(999,32);
				when 35 => sin_data_int <= to_signed(54,32); cos_data_int <= to_signed(998,32);
				when 36 => sin_data_int <= to_signed(55,32); cos_data_int <= to_signed(998,32);
				when 37 => sin_data_int <= to_signed(57,32); cos_data_int <= to_signed(998,32);
				when 38 => sin_data_int <= to_signed(58,32); cos_data_int <= to_signed(998,32);
				when 39 => sin_data_int <= to_signed(60,32); cos_data_int <= to_signed(998,32);
				when 40 => sin_data_int <= to_signed(61,32); cos_data_int <= to_signed(998,32);
				when 41 => sin_data_int <= to_signed(63,32); cos_data_int <= to_signed(998,32);
				when 42 => sin_data_int <= to_signed(64,32); cos_data_int <= to_signed(998,32);
				when 43 => sin_data_int <= to_signed(66,32); cos_data_int <= to_signed(998,32);
				when 44 => sin_data_int <= to_signed(67,32); cos_data_int <= to_signed(998,32);
				when 45 => sin_data_int <= to_signed(69,32); cos_data_int <= to_signed(998,32);
				when 46 => sin_data_int <= to_signed(71,32); cos_data_int <= to_signed(997,32);
				when 47 => sin_data_int <= to_signed(72,32); cos_data_int <= to_signed(997,32);
				when 48 => sin_data_int <= to_signed(74,32); cos_data_int <= to_signed(997,32);
				when 49 => sin_data_int <= to_signed(75,32); cos_data_int <= to_signed(997,32);
				when 50 => sin_data_int <= to_signed(77,32); cos_data_int <= to_signed(997,32);
				when 51 => sin_data_int <= to_signed(78,32); cos_data_int <= to_signed(997,32);
				when 52 => sin_data_int <= to_signed(80,32); cos_data_int <= to_signed(997,32);
				when 53 => sin_data_int <= to_signed(81,32); cos_data_int <= to_signed(997,32);
				when 54 => sin_data_int <= to_signed(83,32); cos_data_int <= to_signed(996,32);
				when 55 => sin_data_int <= to_signed(84,32); cos_data_int <= to_signed(996,32);
				when 56 => sin_data_int <= to_signed(86,32); cos_data_int <= to_signed(996,32);
				when 57 => sin_data_int <= to_signed(87,32); cos_data_int <= to_signed(996,32);
				when 58 => sin_data_int <= to_signed(89,32); cos_data_int <= to_signed(996,32);
				when 59 => sin_data_int <= to_signed(90,32); cos_data_int <= to_signed(996,32);
				when 60 => sin_data_int <= to_signed(92,32); cos_data_int <= to_signed(996,32);
				when 61 => sin_data_int <= to_signed(93,32); cos_data_int <= to_signed(995,32);
				when 62 => sin_data_int <= to_signed(95,32); cos_data_int <= to_signed(995,32);
				when 63 => sin_data_int <= to_signed(96,32); cos_data_int <= to_signed(995,32);
				when 64 => sin_data_int <= to_signed(98,32); cos_data_int <= to_signed(995,32);
				when 65 => sin_data_int <= to_signed(100,32); cos_data_int <= to_signed(995,32);
				when 66 => sin_data_int <= to_signed(101,32); cos_data_int <= to_signed(995,32);
				when 67 => sin_data_int <= to_signed(103,32); cos_data_int <= to_signed(995,32);
				when 68 => sin_data_int <= to_signed(104,32); cos_data_int <= to_signed(994,32);
				when 69 => sin_data_int <= to_signed(106,32); cos_data_int <= to_signed(994,32);
				when 70 => sin_data_int <= to_signed(107,32); cos_data_int <= to_signed(994,32);
				when 71 => sin_data_int <= to_signed(109,32); cos_data_int <= to_signed(994,32);
				when 72 => sin_data_int <= to_signed(110,32); cos_data_int <= to_signed(994,32);
				when 73 => sin_data_int <= to_signed(112,32); cos_data_int <= to_signed(994,32);
				when 74 => sin_data_int <= to_signed(113,32); cos_data_int <= to_signed(993,32);
				when 75 => sin_data_int <= to_signed(115,32); cos_data_int <= to_signed(993,32);
				when 76 => sin_data_int <= to_signed(116,32); cos_data_int <= to_signed(993,32);
				when 77 => sin_data_int <= to_signed(118,32); cos_data_int <= to_signed(993,32);
				when 78 => sin_data_int <= to_signed(119,32); cos_data_int <= to_signed(993,32);
				when 79 => sin_data_int <= to_signed(121,32); cos_data_int <= to_signed(992,32);
				when 80 => sin_data_int <= to_signed(122,32); cos_data_int <= to_signed(992,32);
				when 81 => sin_data_int <= to_signed(124,32); cos_data_int <= to_signed(992,32);
				when 82 => sin_data_int <= to_signed(125,32); cos_data_int <= to_signed(992,32);
				when 83 => sin_data_int <= to_signed(127,32); cos_data_int <= to_signed(992,32);
				when 84 => sin_data_int <= to_signed(128,32); cos_data_int <= to_signed(992,32);
				when 85 => sin_data_int <= to_signed(130,32); cos_data_int <= to_signed(991,32);
				when 86 => sin_data_int <= to_signed(132,32); cos_data_int <= to_signed(991,32);
				when 87 => sin_data_int <= to_signed(133,32); cos_data_int <= to_signed(991,32);
				when 88 => sin_data_int <= to_signed(135,32); cos_data_int <= to_signed(991,32);
				when 89 => sin_data_int <= to_signed(136,32); cos_data_int <= to_signed(990,32);
				when 90 => sin_data_int <= to_signed(138,32); cos_data_int <= to_signed(990,32);
				when 91 => sin_data_int <= to_signed(139,32); cos_data_int <= to_signed(990,32);
				when 92 => sin_data_int <= to_signed(141,32); cos_data_int <= to_signed(990,32);
				when 93 => sin_data_int <= to_signed(142,32); cos_data_int <= to_signed(990,32);
				when 94 => sin_data_int <= to_signed(144,32); cos_data_int <= to_signed(989,32);
				when 95 => sin_data_int <= to_signed(145,32); cos_data_int <= to_signed(989,32);
				when 96 => sin_data_int <= to_signed(147,32); cos_data_int <= to_signed(989,32);
				when 97 => sin_data_int <= to_signed(148,32); cos_data_int <= to_signed(989,32);
				when 98 => sin_data_int <= to_signed(150,32); cos_data_int <= to_signed(988,32);
				when 99 => sin_data_int <= to_signed(151,32); cos_data_int <= to_signed(988,32);
				when 100 => sin_data_int <= to_signed(153,32); cos_data_int <= to_signed(988,32);
				when 101 => sin_data_int <= to_signed(154,32); cos_data_int <= to_signed(988,32);
				when 102 => sin_data_int <= to_signed(156,32); cos_data_int <= to_signed(988,32);
				when 103 => sin_data_int <= to_signed(157,32); cos_data_int <= to_signed(987,32);
				when 104 => sin_data_int <= to_signed(159,32); cos_data_int <= to_signed(987,32);
				when 105 => sin_data_int <= to_signed(160,32); cos_data_int <= to_signed(987,32);
				when 106 => sin_data_int <= to_signed(162,32); cos_data_int <= to_signed(987,32);
				when 107 => sin_data_int <= to_signed(163,32); cos_data_int <= to_signed(986,32);
				when 108 => sin_data_int <= to_signed(165,32); cos_data_int <= to_signed(986,32);
				when 109 => sin_data_int <= to_signed(166,32); cos_data_int <= to_signed(986,32);
				when 110 => sin_data_int <= to_signed(168,32); cos_data_int <= to_signed(986,32);
				when 111 => sin_data_int <= to_signed(169,32); cos_data_int <= to_signed(985,32);
				when 112 => sin_data_int <= to_signed(171,32); cos_data_int <= to_signed(985,32);
				when 113 => sin_data_int <= to_signed(172,32); cos_data_int <= to_signed(985,32);
				when 114 => sin_data_int <= to_signed(174,32); cos_data_int <= to_signed(984,32);
				when 115 => sin_data_int <= to_signed(175,32); cos_data_int <= to_signed(984,32);
				when 116 => sin_data_int <= to_signed(177,32); cos_data_int <= to_signed(984,32);
				when 117 => sin_data_int <= to_signed(179,32); cos_data_int <= to_signed(984,32);
				when 118 => sin_data_int <= to_signed(180,32); cos_data_int <= to_signed(983,32);
				when 119 => sin_data_int <= to_signed(182,32); cos_data_int <= to_signed(983,32);
				when 120 => sin_data_int <= to_signed(183,32); cos_data_int <= to_signed(983,32);
				when 121 => sin_data_int <= to_signed(185,32); cos_data_int <= to_signed(983,32);
				when 122 => sin_data_int <= to_signed(186,32); cos_data_int <= to_signed(982,32);
				when 123 => sin_data_int <= to_signed(188,32); cos_data_int <= to_signed(982,32);
				when 124 => sin_data_int <= to_signed(189,32); cos_data_int <= to_signed(982,32);
				when 125 => sin_data_int <= to_signed(191,32); cos_data_int <= to_signed(981,32);
				when 126 => sin_data_int <= to_signed(192,32); cos_data_int <= to_signed(981,32);
				when 127 => sin_data_int <= to_signed(194,32); cos_data_int <= to_signed(981,32);
				when 128 => sin_data_int <= to_signed(195,32); cos_data_int <= to_signed(980,32);
				when 129 => sin_data_int <= to_signed(197,32); cos_data_int <= to_signed(980,32);
				when 130 => sin_data_int <= to_signed(198,32); cos_data_int <= to_signed(980,32);
				when 131 => sin_data_int <= to_signed(200,32); cos_data_int <= to_signed(980,32);
				when 132 => sin_data_int <= to_signed(201,32); cos_data_int <= to_signed(979,32);
				when 133 => sin_data_int <= to_signed(203,32); cos_data_int <= to_signed(979,32);
				when 134 => sin_data_int <= to_signed(204,32); cos_data_int <= to_signed(979,32);
				when 135 => sin_data_int <= to_signed(206,32); cos_data_int <= to_signed(978,32);
				when 136 => sin_data_int <= to_signed(207,32); cos_data_int <= to_signed(978,32);
				when 137 => sin_data_int <= to_signed(209,32); cos_data_int <= to_signed(978,32);
				when 138 => sin_data_int <= to_signed(210,32); cos_data_int <= to_signed(977,32);
				when 139 => sin_data_int <= to_signed(212,32); cos_data_int <= to_signed(977,32);
				when 140 => sin_data_int <= to_signed(213,32); cos_data_int <= to_signed(977,32);
				when 141 => sin_data_int <= to_signed(215,32); cos_data_int <= to_signed(976,32);
				when 142 => sin_data_int <= to_signed(216,32); cos_data_int <= to_signed(976,32);
				when 143 => sin_data_int <= to_signed(218,32); cos_data_int <= to_signed(976,32);
				when 144 => sin_data_int <= to_signed(219,32); cos_data_int <= to_signed(975,32);
				when 145 => sin_data_int <= to_signed(221,32); cos_data_int <= to_signed(975,32);
				when 146 => sin_data_int <= to_signed(222,32); cos_data_int <= to_signed(975,32);
				when 147 => sin_data_int <= to_signed(224,32); cos_data_int <= to_signed(974,32);
				when 148 => sin_data_int <= to_signed(225,32); cos_data_int <= to_signed(974,32);
				when 149 => sin_data_int <= to_signed(227,32); cos_data_int <= to_signed(974,32);
				when 150 => sin_data_int <= to_signed(228,32); cos_data_int <= to_signed(973,32);
				when 151 => sin_data_int <= to_signed(230,32); cos_data_int <= to_signed(973,32);
				when 152 => sin_data_int <= to_signed(231,32); cos_data_int <= to_signed(973,32);
				when 153 => sin_data_int <= to_signed(233,32); cos_data_int <= to_signed(972,32);
				when 154 => sin_data_int <= to_signed(234,32); cos_data_int <= to_signed(972,32);
				when 155 => sin_data_int <= to_signed(236,32); cos_data_int <= to_signed(972,32);
				when 156 => sin_data_int <= to_signed(237,32); cos_data_int <= to_signed(971,32);
				when 157 => sin_data_int <= to_signed(239,32); cos_data_int <= to_signed(971,32);
				when 158 => sin_data_int <= to_signed(240,32); cos_data_int <= to_signed(970,32);
				when 159 => sin_data_int <= to_signed(241,32); cos_data_int <= to_signed(970,32);
				when 160 => sin_data_int <= to_signed(243,32); cos_data_int <= to_signed(970,32);
				when 161 => sin_data_int <= to_signed(244,32); cos_data_int <= to_signed(969,32);
				when 162 => sin_data_int <= to_signed(246,32); cos_data_int <= to_signed(969,32);
				when 163 => sin_data_int <= to_signed(247,32); cos_data_int <= to_signed(969,32);
				when 164 => sin_data_int <= to_signed(249,32); cos_data_int <= to_signed(968,32);
				when 165 => sin_data_int <= to_signed(250,32); cos_data_int <= to_signed(968,32);
				when 166 => sin_data_int <= to_signed(252,32); cos_data_int <= to_signed(967,32);
				when 167 => sin_data_int <= to_signed(253,32); cos_data_int <= to_signed(967,32);
				when 168 => sin_data_int <= to_signed(255,32); cos_data_int <= to_signed(967,32);
				when 169 => sin_data_int <= to_signed(256,32); cos_data_int <= to_signed(966,32);
				when 170 => sin_data_int <= to_signed(258,32); cos_data_int <= to_signed(966,32);
				when 171 => sin_data_int <= to_signed(259,32); cos_data_int <= to_signed(965,32);
				when 172 => sin_data_int <= to_signed(261,32); cos_data_int <= to_signed(965,32);
				when 173 => sin_data_int <= to_signed(262,32); cos_data_int <= to_signed(965,32);
				when 174 => sin_data_int <= to_signed(264,32); cos_data_int <= to_signed(964,32);
				when 175 => sin_data_int <= to_signed(265,32); cos_data_int <= to_signed(964,32);
				when 176 => sin_data_int <= to_signed(267,32); cos_data_int <= to_signed(963,32);
				when 177 => sin_data_int <= to_signed(268,32); cos_data_int <= to_signed(963,32);
				when 178 => sin_data_int <= to_signed(270,32); cos_data_int <= to_signed(963,32);
				when 179 => sin_data_int <= to_signed(271,32); cos_data_int <= to_signed(962,32);
				when 180 => sin_data_int <= to_signed(273,32); cos_data_int <= to_signed(962,32);
				when 181 => sin_data_int <= to_signed(274,32); cos_data_int <= to_signed(961,32);
				when 182 => sin_data_int <= to_signed(276,32); cos_data_int <= to_signed(961,32);
				when 183 => sin_data_int <= to_signed(277,32); cos_data_int <= to_signed(960,32);
				when 184 => sin_data_int <= to_signed(279,32); cos_data_int <= to_signed(960,32);
				when 185 => sin_data_int <= to_signed(280,32); cos_data_int <= to_signed(960,32);
				when 186 => sin_data_int <= to_signed(281,32); cos_data_int <= to_signed(959,32);
				when 187 => sin_data_int <= to_signed(283,32); cos_data_int <= to_signed(959,32);
				when 188 => sin_data_int <= to_signed(284,32); cos_data_int <= to_signed(958,32);
				when 189 => sin_data_int <= to_signed(286,32); cos_data_int <= to_signed(958,32);
				when 190 => sin_data_int <= to_signed(287,32); cos_data_int <= to_signed(957,32);
				when 191 => sin_data_int <= to_signed(289,32); cos_data_int <= to_signed(957,32);
				when 192 => sin_data_int <= to_signed(290,32); cos_data_int <= to_signed(956,32);
				when 193 => sin_data_int <= to_signed(292,32); cos_data_int <= to_signed(956,32);
				when 194 => sin_data_int <= to_signed(293,32); cos_data_int <= to_signed(956,32);
				when 195 => sin_data_int <= to_signed(295,32); cos_data_int <= to_signed(955,32);
				when 196 => sin_data_int <= to_signed(296,32); cos_data_int <= to_signed(955,32);
				when 197 => sin_data_int <= to_signed(298,32); cos_data_int <= to_signed(954,32);
				when 198 => sin_data_int <= to_signed(299,32); cos_data_int <= to_signed(954,32);
				when 199 => sin_data_int <= to_signed(301,32); cos_data_int <= to_signed(953,32);
				when 200 => sin_data_int <= to_signed(302,32); cos_data_int <= to_signed(953,32);
				when 201 => sin_data_int <= to_signed(303,32); cos_data_int <= to_signed(952,32);
				when 202 => sin_data_int <= to_signed(305,32); cos_data_int <= to_signed(952,32);
				when 203 => sin_data_int <= to_signed(306,32); cos_data_int <= to_signed(951,32);
				when 204 => sin_data_int <= to_signed(308,32); cos_data_int <= to_signed(951,32);
				when 205 => sin_data_int <= to_signed(309,32); cos_data_int <= to_signed(950,32);
				when 206 => sin_data_int <= to_signed(311,32); cos_data_int <= to_signed(950,32);
				when 207 => sin_data_int <= to_signed(312,32); cos_data_int <= to_signed(950,32);
				when 208 => sin_data_int <= to_signed(314,32); cos_data_int <= to_signed(949,32);
				when 209 => sin_data_int <= to_signed(315,32); cos_data_int <= to_signed(949,32);
				when 210 => sin_data_int <= to_signed(317,32); cos_data_int <= to_signed(948,32);
				when 211 => sin_data_int <= to_signed(318,32); cos_data_int <= to_signed(948,32);
				when 212 => sin_data_int <= to_signed(320,32); cos_data_int <= to_signed(947,32);
				when 213 => sin_data_int <= to_signed(321,32); cos_data_int <= to_signed(947,32);
				when 214 => sin_data_int <= to_signed(322,32); cos_data_int <= to_signed(946,32);
				when 215 => sin_data_int <= to_signed(324,32); cos_data_int <= to_signed(946,32);
				when 216 => sin_data_int <= to_signed(325,32); cos_data_int <= to_signed(945,32);
				when 217 => sin_data_int <= to_signed(327,32); cos_data_int <= to_signed(945,32);
				when 218 => sin_data_int <= to_signed(328,32); cos_data_int <= to_signed(944,32);
				when 219 => sin_data_int <= to_signed(330,32); cos_data_int <= to_signed(944,32);
				when 220 => sin_data_int <= to_signed(331,32); cos_data_int <= to_signed(943,32);
				when 221 => sin_data_int <= to_signed(333,32); cos_data_int <= to_signed(943,32);
				when 222 => sin_data_int <= to_signed(334,32); cos_data_int <= to_signed(942,32);
				when 223 => sin_data_int <= to_signed(335,32); cos_data_int <= to_signed(942,32);
				when 224 => sin_data_int <= to_signed(337,32); cos_data_int <= to_signed(941,32);
				when 225 => sin_data_int <= to_signed(338,32); cos_data_int <= to_signed(941,32);
				when 226 => sin_data_int <= to_signed(340,32); cos_data_int <= to_signed(940,32);
				when 227 => sin_data_int <= to_signed(341,32); cos_data_int <= to_signed(939,32);
				when 228 => sin_data_int <= to_signed(343,32); cos_data_int <= to_signed(939,32);
				when 229 => sin_data_int <= to_signed(344,32); cos_data_int <= to_signed(938,32);
				when 230 => sin_data_int <= to_signed(346,32); cos_data_int <= to_signed(938,32);
				when 231 => sin_data_int <= to_signed(347,32); cos_data_int <= to_signed(937,32);
				when 232 => sin_data_int <= to_signed(348,32); cos_data_int <= to_signed(937,32);
				when 233 => sin_data_int <= to_signed(350,32); cos_data_int <= to_signed(936,32);
				when 234 => sin_data_int <= to_signed(351,32); cos_data_int <= to_signed(936,32);
				when 235 => sin_data_int <= to_signed(353,32); cos_data_int <= to_signed(935,32);
				when 236 => sin_data_int <= to_signed(354,32); cos_data_int <= to_signed(935,32);
				when 237 => sin_data_int <= to_signed(356,32); cos_data_int <= to_signed(934,32);
				when 238 => sin_data_int <= to_signed(357,32); cos_data_int <= to_signed(934,32);
				when 239 => sin_data_int <= to_signed(358,32); cos_data_int <= to_signed(933,32);
				when 240 => sin_data_int <= to_signed(360,32); cos_data_int <= to_signed(932,32);
				when 241 => sin_data_int <= to_signed(361,32); cos_data_int <= to_signed(932,32);
				when 242 => sin_data_int <= to_signed(363,32); cos_data_int <= to_signed(931,32);
				when 243 => sin_data_int <= to_signed(364,32); cos_data_int <= to_signed(931,32);
				when 244 => sin_data_int <= to_signed(366,32); cos_data_int <= to_signed(930,32);
				when 245 => sin_data_int <= to_signed(367,32); cos_data_int <= to_signed(930,32);
				when 246 => sin_data_int <= to_signed(368,32); cos_data_int <= to_signed(929,32);
				when 247 => sin_data_int <= to_signed(370,32); cos_data_int <= to_signed(929,32);
				when 248 => sin_data_int <= to_signed(371,32); cos_data_int <= to_signed(928,32);
				when 249 => sin_data_int <= to_signed(373,32); cos_data_int <= to_signed(927,32);
				when 250 => sin_data_int <= to_signed(374,32); cos_data_int <= to_signed(927,32);
				when 251 => sin_data_int <= to_signed(376,32); cos_data_int <= to_signed(926,32);
				when 252 => sin_data_int <= to_signed(377,32); cos_data_int <= to_signed(926,32);
				when 253 => sin_data_int <= to_signed(378,32); cos_data_int <= to_signed(925,32);
				when 254 => sin_data_int <= to_signed(380,32); cos_data_int <= to_signed(924,32);
				when 255 => sin_data_int <= to_signed(381,32); cos_data_int <= to_signed(924,32);
				when 256 => sin_data_int <= to_signed(383,32); cos_data_int <= to_signed(923,32);
				when 257 => sin_data_int <= to_signed(384,32); cos_data_int <= to_signed(923,32);
				when 258 => sin_data_int <= to_signed(386,32); cos_data_int <= to_signed(922,32);
				when 259 => sin_data_int <= to_signed(387,32); cos_data_int <= to_signed(922,32);
				when 260 => sin_data_int <= to_signed(388,32); cos_data_int <= to_signed(921,32);
				when 261 => sin_data_int <= to_signed(390,32); cos_data_int <= to_signed(920,32);
				when 262 => sin_data_int <= to_signed(391,32); cos_data_int <= to_signed(920,32);
				when 263 => sin_data_int <= to_signed(393,32); cos_data_int <= to_signed(919,32);
				when 264 => sin_data_int <= to_signed(394,32); cos_data_int <= to_signed(919,32);
				when 265 => sin_data_int <= to_signed(395,32); cos_data_int <= to_signed(918,32);
				when 266 => sin_data_int <= to_signed(397,32); cos_data_int <= to_signed(917,32);
				when 267 => sin_data_int <= to_signed(398,32); cos_data_int <= to_signed(917,32);
				when 268 => sin_data_int <= to_signed(400,32); cos_data_int <= to_signed(916,32);
				when 269 => sin_data_int <= to_signed(401,32); cos_data_int <= to_signed(915,32);
				when 270 => sin_data_int <= to_signed(402,32); cos_data_int <= to_signed(915,32);
				when 271 => sin_data_int <= to_signed(404,32); cos_data_int <= to_signed(914,32);
				when 272 => sin_data_int <= to_signed(405,32); cos_data_int <= to_signed(914,32);
				when 273 => sin_data_int <= to_signed(407,32); cos_data_int <= to_signed(913,32);
				when 274 => sin_data_int <= to_signed(408,32); cos_data_int <= to_signed(912,32);
				when 275 => sin_data_int <= to_signed(409,32); cos_data_int <= to_signed(912,32);
				when 276 => sin_data_int <= to_signed(411,32); cos_data_int <= to_signed(911,32);
				when 277 => sin_data_int <= to_signed(412,32); cos_data_int <= to_signed(910,32);
				when 278 => sin_data_int <= to_signed(414,32); cos_data_int <= to_signed(910,32);
				when 279 => sin_data_int <= to_signed(415,32); cos_data_int <= to_signed(909,32);
				when 280 => sin_data_int <= to_signed(416,32); cos_data_int <= to_signed(909,32);
				when 281 => sin_data_int <= to_signed(418,32); cos_data_int <= to_signed(908,32);
				when 282 => sin_data_int <= to_signed(419,32); cos_data_int <= to_signed(907,32);
				when 283 => sin_data_int <= to_signed(421,32); cos_data_int <= to_signed(907,32);
				when 284 => sin_data_int <= to_signed(422,32); cos_data_int <= to_signed(906,32);
				when 285 => sin_data_int <= to_signed(423,32); cos_data_int <= to_signed(905,32);
				when 286 => sin_data_int <= to_signed(425,32); cos_data_int <= to_signed(905,32);
				when 287 => sin_data_int <= to_signed(426,32); cos_data_int <= to_signed(904,32);
				when 288 => sin_data_int <= to_signed(428,32); cos_data_int <= to_signed(903,32);
				when 289 => sin_data_int <= to_signed(429,32); cos_data_int <= to_signed(903,32);
				when 290 => sin_data_int <= to_signed(430,32); cos_data_int <= to_signed(902,32);
				when 291 => sin_data_int <= to_signed(432,32); cos_data_int <= to_signed(901,32);
				when 292 => sin_data_int <= to_signed(433,32); cos_data_int <= to_signed(901,32);
				when 293 => sin_data_int <= to_signed(434,32); cos_data_int <= to_signed(900,32);
				when 294 => sin_data_int <= to_signed(436,32); cos_data_int <= to_signed(899,32);
				when 295 => sin_data_int <= to_signed(437,32); cos_data_int <= to_signed(899,32);
				when 296 => sin_data_int <= to_signed(439,32); cos_data_int <= to_signed(898,32);
				when 297 => sin_data_int <= to_signed(440,32); cos_data_int <= to_signed(897,32);
				when 298 => sin_data_int <= to_signed(441,32); cos_data_int <= to_signed(897,32);
				when 299 => sin_data_int <= to_signed(443,32); cos_data_int <= to_signed(896,32);
				when 300 => sin_data_int <= to_signed(444,32); cos_data_int <= to_signed(895,32);
				when 301 => sin_data_int <= to_signed(445,32); cos_data_int <= to_signed(895,32);
				when 302 => sin_data_int <= to_signed(447,32); cos_data_int <= to_signed(894,32);
				when 303 => sin_data_int <= to_signed(448,32); cos_data_int <= to_signed(893,32);
				when 304 => sin_data_int <= to_signed(450,32); cos_data_int <= to_signed(893,32);
				when 305 => sin_data_int <= to_signed(451,32); cos_data_int <= to_signed(892,32);
				when 306 => sin_data_int <= to_signed(452,32); cos_data_int <= to_signed(891,32);
				when 307 => sin_data_int <= to_signed(454,32); cos_data_int <= to_signed(890,32);
				when 308 => sin_data_int <= to_signed(455,32); cos_data_int <= to_signed(890,32);
				when 309 => sin_data_int <= to_signed(456,32); cos_data_int <= to_signed(889,32);
				when 310 => sin_data_int <= to_signed(458,32); cos_data_int <= to_signed(888,32);
				when 311 => sin_data_int <= to_signed(459,32); cos_data_int <= to_signed(888,32);
				when 312 => sin_data_int <= to_signed(461,32); cos_data_int <= to_signed(887,32);
				when 313 => sin_data_int <= to_signed(462,32); cos_data_int <= to_signed(886,32);
				when 314 => sin_data_int <= to_signed(463,32); cos_data_int <= to_signed(886,32);
				when 315 => sin_data_int <= to_signed(465,32); cos_data_int <= to_signed(885,32);
				when 316 => sin_data_int <= to_signed(466,32); cos_data_int <= to_signed(884,32);
				when 317 => sin_data_int <= to_signed(467,32); cos_data_int <= to_signed(883,32);
				when 318 => sin_data_int <= to_signed(469,32); cos_data_int <= to_signed(883,32);
				when 319 => sin_data_int <= to_signed(470,32); cos_data_int <= to_signed(882,32);
				when 320 => sin_data_int <= to_signed(471,32); cos_data_int <= to_signed(881,32);
				when 321 => sin_data_int <= to_signed(473,32); cos_data_int <= to_signed(880,32);
				when 322 => sin_data_int <= to_signed(474,32); cos_data_int <= to_signed(880,32);
				when 323 => sin_data_int <= to_signed(475,32); cos_data_int <= to_signed(879,32);
				when 324 => sin_data_int <= to_signed(477,32); cos_data_int <= to_signed(878,32);
				when 325 => sin_data_int <= to_signed(478,32); cos_data_int <= to_signed(878,32);
				when 326 => sin_data_int <= to_signed(479,32); cos_data_int <= to_signed(877,32);
				when 327 => sin_data_int <= to_signed(481,32); cos_data_int <= to_signed(876,32);
				when 328 => sin_data_int <= to_signed(482,32); cos_data_int <= to_signed(875,32);
				when 329 => sin_data_int <= to_signed(484,32); cos_data_int <= to_signed(875,32);
				when 330 => sin_data_int <= to_signed(485,32); cos_data_int <= to_signed(874,32);
				when 331 => sin_data_int <= to_signed(486,32); cos_data_int <= to_signed(873,32);
				when 332 => sin_data_int <= to_signed(488,32); cos_data_int <= to_signed(872,32);
				when 333 => sin_data_int <= to_signed(489,32); cos_data_int <= to_signed(872,32);
				when 334 => sin_data_int <= to_signed(490,32); cos_data_int <= to_signed(871,32);
				when 335 => sin_data_int <= to_signed(492,32); cos_data_int <= to_signed(870,32);
				when 336 => sin_data_int <= to_signed(493,32); cos_data_int <= to_signed(869,32);
				when 337 => sin_data_int <= to_signed(494,32); cos_data_int <= to_signed(869,32);
				when 338 => sin_data_int <= to_signed(496,32); cos_data_int <= to_signed(868,32);
				when 339 => sin_data_int <= to_signed(497,32); cos_data_int <= to_signed(867,32);
				when 340 => sin_data_int <= to_signed(498,32); cos_data_int <= to_signed(866,32);
				when 341 => sin_data_int <= to_signed(500,32); cos_data_int <= to_signed(866,32);
				when 342 => sin_data_int <= to_signed(501,32); cos_data_int <= to_signed(865,32);
				when 343 => sin_data_int <= to_signed(502,32); cos_data_int <= to_signed(864,32);
				when 344 => sin_data_int <= to_signed(504,32); cos_data_int <= to_signed(863,32);
				when 345 => sin_data_int <= to_signed(505,32); cos_data_int <= to_signed(862,32);
				when 346 => sin_data_int <= to_signed(506,32); cos_data_int <= to_signed(862,32);
				when 347 => sin_data_int <= to_signed(508,32); cos_data_int <= to_signed(861,32);
				when 348 => sin_data_int <= to_signed(509,32); cos_data_int <= to_signed(860,32);
				when 349 => sin_data_int <= to_signed(510,32); cos_data_int <= to_signed(859,32);
				when 350 => sin_data_int <= to_signed(511,32); cos_data_int <= to_signed(859,32);
				when 351 => sin_data_int <= to_signed(513,32); cos_data_int <= to_signed(858,32);
				when 352 => sin_data_int <= to_signed(514,32); cos_data_int <= to_signed(857,32);
				when 353 => sin_data_int <= to_signed(515,32); cos_data_int <= to_signed(856,32);
				when 354 => sin_data_int <= to_signed(517,32); cos_data_int <= to_signed(855,32);
				when 355 => sin_data_int <= to_signed(518,32); cos_data_int <= to_signed(855,32);
				when 356 => sin_data_int <= to_signed(519,32); cos_data_int <= to_signed(854,32);
				when 357 => sin_data_int <= to_signed(521,32); cos_data_int <= to_signed(853,32);
				when 358 => sin_data_int <= to_signed(522,32); cos_data_int <= to_signed(852,32);
				when 359 => sin_data_int <= to_signed(523,32); cos_data_int <= to_signed(851,32);
				when 360 => sin_data_int <= to_signed(525,32); cos_data_int <= to_signed(851,32);
				when 361 => sin_data_int <= to_signed(526,32); cos_data_int <= to_signed(850,32);
				when 362 => sin_data_int <= to_signed(527,32); cos_data_int <= to_signed(849,32);
				when 363 => sin_data_int <= to_signed(529,32); cos_data_int <= to_signed(848,32);
				when 364 => sin_data_int <= to_signed(530,32); cos_data_int <= to_signed(847,32);
				when 365 => sin_data_int <= to_signed(531,32); cos_data_int <= to_signed(846,32);
				when 366 => sin_data_int <= to_signed(532,32); cos_data_int <= to_signed(846,32);
				when 367 => sin_data_int <= to_signed(534,32); cos_data_int <= to_signed(845,32);
				when 368 => sin_data_int <= to_signed(535,32); cos_data_int <= to_signed(844,32);
				when 369 => sin_data_int <= to_signed(536,32); cos_data_int <= to_signed(843,32);
				when 370 => sin_data_int <= to_signed(538,32); cos_data_int <= to_signed(842,32);
				when 371 => sin_data_int <= to_signed(539,32); cos_data_int <= to_signed(842,32);
				when 372 => sin_data_int <= to_signed(540,32); cos_data_int <= to_signed(841,32);
				when 373 => sin_data_int <= to_signed(541,32); cos_data_int <= to_signed(840,32);
				when 374 => sin_data_int <= to_signed(543,32); cos_data_int <= to_signed(839,32);
				when 375 => sin_data_int <= to_signed(544,32); cos_data_int <= to_signed(838,32);
				when 376 => sin_data_int <= to_signed(545,32); cos_data_int <= to_signed(837,32);
				when 377 => sin_data_int <= to_signed(547,32); cos_data_int <= to_signed(837,32);
				when 378 => sin_data_int <= to_signed(548,32); cos_data_int <= to_signed(836,32);
				when 379 => sin_data_int <= to_signed(549,32); cos_data_int <= to_signed(835,32);
				when 380 => sin_data_int <= to_signed(550,32); cos_data_int <= to_signed(834,32);
				when 381 => sin_data_int <= to_signed(552,32); cos_data_int <= to_signed(833,32);
				when 382 => sin_data_int <= to_signed(553,32); cos_data_int <= to_signed(832,32);
				when 383 => sin_data_int <= to_signed(554,32); cos_data_int <= to_signed(831,32);
				when 384 => sin_data_int <= to_signed(556,32); cos_data_int <= to_signed(831,32);
				when 385 => sin_data_int <= to_signed(557,32); cos_data_int <= to_signed(830,32);
				when 386 => sin_data_int <= to_signed(558,32); cos_data_int <= to_signed(829,32);
				when 387 => sin_data_int <= to_signed(559,32); cos_data_int <= to_signed(828,32);
				when 388 => sin_data_int <= to_signed(561,32); cos_data_int <= to_signed(827,32);
				when 389 => sin_data_int <= to_signed(562,32); cos_data_int <= to_signed(826,32);
				when 390 => sin_data_int <= to_signed(563,32); cos_data_int <= to_signed(825,32);
				when 391 => sin_data_int <= to_signed(564,32); cos_data_int <= to_signed(825,32);
				when 392 => sin_data_int <= to_signed(566,32); cos_data_int <= to_signed(824,32);
				when 393 => sin_data_int <= to_signed(567,32); cos_data_int <= to_signed(823,32);
				when 394 => sin_data_int <= to_signed(568,32); cos_data_int <= to_signed(822,32);
				when 395 => sin_data_int <= to_signed(570,32); cos_data_int <= to_signed(821,32);
				when 396 => sin_data_int <= to_signed(571,32); cos_data_int <= to_signed(820,32);
				when 397 => sin_data_int <= to_signed(572,32); cos_data_int <= to_signed(819,32);
				when 398 => sin_data_int <= to_signed(573,32); cos_data_int <= to_signed(818,32);
				when 399 => sin_data_int <= to_signed(575,32); cos_data_int <= to_signed(818,32);
				when 400 => sin_data_int <= to_signed(576,32); cos_data_int <= to_signed(817,32);
				when 401 => sin_data_int <= to_signed(577,32); cos_data_int <= to_signed(816,32);
				when 402 => sin_data_int <= to_signed(578,32); cos_data_int <= to_signed(815,32);
				when 403 => sin_data_int <= to_signed(580,32); cos_data_int <= to_signed(814,32);
				when 404 => sin_data_int <= to_signed(581,32); cos_data_int <= to_signed(813,32);
				when 405 => sin_data_int <= to_signed(582,32); cos_data_int <= to_signed(812,32);
				when 406 => sin_data_int <= to_signed(583,32); cos_data_int <= to_signed(811,32);
				when 407 => sin_data_int <= to_signed(585,32); cos_data_int <= to_signed(810,32);
				when 408 => sin_data_int <= to_signed(586,32); cos_data_int <= to_signed(810,32);
				when 409 => sin_data_int <= to_signed(587,32); cos_data_int <= to_signed(809,32);
				when 410 => sin_data_int <= to_signed(588,32); cos_data_int <= to_signed(808,32);
				when 411 => sin_data_int <= to_signed(590,32); cos_data_int <= to_signed(807,32);
				when 412 => sin_data_int <= to_signed(591,32); cos_data_int <= to_signed(806,32);
				when 413 => sin_data_int <= to_signed(592,32); cos_data_int <= to_signed(805,32);
				when 414 => sin_data_int <= to_signed(593,32); cos_data_int <= to_signed(804,32);
				when 415 => sin_data_int <= to_signed(594,32); cos_data_int <= to_signed(803,32);
				when 416 => sin_data_int <= to_signed(596,32); cos_data_int <= to_signed(802,32);
				when 417 => sin_data_int <= to_signed(597,32); cos_data_int <= to_signed(801,32);
				when 418 => sin_data_int <= to_signed(598,32); cos_data_int <= to_signed(800,32);
				when 419 => sin_data_int <= to_signed(599,32); cos_data_int <= to_signed(800,32);
				when 420 => sin_data_int <= to_signed(601,32); cos_data_int <= to_signed(799,32);
				when 421 => sin_data_int <= to_signed(602,32); cos_data_int <= to_signed(798,32);
				when 422 => sin_data_int <= to_signed(603,32); cos_data_int <= to_signed(797,32);
				when 423 => sin_data_int <= to_signed(604,32); cos_data_int <= to_signed(796,32);
				when 424 => sin_data_int <= to_signed(606,32); cos_data_int <= to_signed(795,32);
				when 425 => sin_data_int <= to_signed(607,32); cos_data_int <= to_signed(794,32);
				when 426 => sin_data_int <= to_signed(608,32); cos_data_int <= to_signed(793,32);
				when 427 => sin_data_int <= to_signed(609,32); cos_data_int <= to_signed(792,32);
				when 428 => sin_data_int <= to_signed(610,32); cos_data_int <= to_signed(791,32);
				when 429 => sin_data_int <= to_signed(612,32); cos_data_int <= to_signed(790,32);
				when 430 => sin_data_int <= to_signed(613,32); cos_data_int <= to_signed(789,32);
				when 431 => sin_data_int <= to_signed(614,32); cos_data_int <= to_signed(788,32);
				when 432 => sin_data_int <= to_signed(615,32); cos_data_int <= to_signed(787,32);
				when 433 => sin_data_int <= to_signed(616,32); cos_data_int <= to_signed(786,32);
				when 434 => sin_data_int <= to_signed(618,32); cos_data_int <= to_signed(786,32);
				when 435 => sin_data_int <= to_signed(619,32); cos_data_int <= to_signed(785,32);
				when 436 => sin_data_int <= to_signed(620,32); cos_data_int <= to_signed(784,32);
				when 437 => sin_data_int <= to_signed(621,32); cos_data_int <= to_signed(783,32);
				when 438 => sin_data_int <= to_signed(622,32); cos_data_int <= to_signed(782,32);
				when 439 => sin_data_int <= to_signed(624,32); cos_data_int <= to_signed(781,32);
				when 440 => sin_data_int <= to_signed(625,32); cos_data_int <= to_signed(780,32);
				when 441 => sin_data_int <= to_signed(626,32); cos_data_int <= to_signed(779,32);
				when 442 => sin_data_int <= to_signed(627,32); cos_data_int <= to_signed(778,32);
				when 443 => sin_data_int <= to_signed(628,32); cos_data_int <= to_signed(777,32);
				when 444 => sin_data_int <= to_signed(630,32); cos_data_int <= to_signed(776,32);
				when 445 => sin_data_int <= to_signed(631,32); cos_data_int <= to_signed(775,32);
				when 446 => sin_data_int <= to_signed(632,32); cos_data_int <= to_signed(774,32);
				when 447 => sin_data_int <= to_signed(633,32); cos_data_int <= to_signed(773,32);
				when 448 => sin_data_int <= to_signed(634,32); cos_data_int <= to_signed(772,32);
				when 449 => sin_data_int <= to_signed(636,32); cos_data_int <= to_signed(771,32);
				when 450 => sin_data_int <= to_signed(637,32); cos_data_int <= to_signed(770,32);
				when 451 => sin_data_int <= to_signed(638,32); cos_data_int <= to_signed(769,32);
				when 452 => sin_data_int <= to_signed(639,32); cos_data_int <= to_signed(768,32);
				when 453 => sin_data_int <= to_signed(640,32); cos_data_int <= to_signed(767,32);
				when 454 => sin_data_int <= to_signed(641,32); cos_data_int <= to_signed(766,32);
				when 455 => sin_data_int <= to_signed(643,32); cos_data_int <= to_signed(765,32);
				when 456 => sin_data_int <= to_signed(644,32); cos_data_int <= to_signed(764,32);
				when 457 => sin_data_int <= to_signed(645,32); cos_data_int <= to_signed(763,32);
				when 458 => sin_data_int <= to_signed(646,32); cos_data_int <= to_signed(762,32);
				when 459 => sin_data_int <= to_signed(647,32); cos_data_int <= to_signed(761,32);
				when 460 => sin_data_int <= to_signed(649,32); cos_data_int <= to_signed(760,32);
				when 461 => sin_data_int <= to_signed(650,32); cos_data_int <= to_signed(759,32);
				when 462 => sin_data_int <= to_signed(651,32); cos_data_int <= to_signed(758,32);
				when 463 => sin_data_int <= to_signed(652,32); cos_data_int <= to_signed(757,32);
				when 464 => sin_data_int <= to_signed(653,32); cos_data_int <= to_signed(756,32);
				when 465 => sin_data_int <= to_signed(654,32); cos_data_int <= to_signed(755,32);
				when 466 => sin_data_int <= to_signed(655,32); cos_data_int <= to_signed(754,32);
				when 467 => sin_data_int <= to_signed(657,32); cos_data_int <= to_signed(753,32);
				when 468 => sin_data_int <= to_signed(658,32); cos_data_int <= to_signed(752,32);
				when 469 => sin_data_int <= to_signed(659,32); cos_data_int <= to_signed(751,32);
				when 470 => sin_data_int <= to_signed(660,32); cos_data_int <= to_signed(750,32);
				when 471 => sin_data_int <= to_signed(661,32); cos_data_int <= to_signed(749,32);
				when 472 => sin_data_int <= to_signed(662,32); cos_data_int <= to_signed(748,32);
				when 473 => sin_data_int <= to_signed(664,32); cos_data_int <= to_signed(747,32);
				when 474 => sin_data_int <= to_signed(665,32); cos_data_int <= to_signed(746,32);
				when 475 => sin_data_int <= to_signed(666,32); cos_data_int <= to_signed(745,32);
				when 476 => sin_data_int <= to_signed(667,32); cos_data_int <= to_signed(744,32);
				when 477 => sin_data_int <= to_signed(668,32); cos_data_int <= to_signed(743,32);
				when 478 => sin_data_int <= to_signed(669,32); cos_data_int <= to_signed(742,32);
				when 479 => sin_data_int <= to_signed(670,32); cos_data_int <= to_signed(741,32);
				when 480 => sin_data_int <= to_signed(672,32); cos_data_int <= to_signed(740,32);
				when 481 => sin_data_int <= to_signed(673,32); cos_data_int <= to_signed(739,32);
				when 482 => sin_data_int <= to_signed(674,32); cos_data_int <= to_signed(738,32);
				when 483 => sin_data_int <= to_signed(675,32); cos_data_int <= to_signed(737,32);
				when 484 => sin_data_int <= to_signed(676,32); cos_data_int <= to_signed(736,32);
				when 485 => sin_data_int <= to_signed(677,32); cos_data_int <= to_signed(735,32);
				when 486 => sin_data_int <= to_signed(678,32); cos_data_int <= to_signed(734,32);
				when 487 => sin_data_int <= to_signed(679,32); cos_data_int <= to_signed(733,32);
				when 488 => sin_data_int <= to_signed(681,32); cos_data_int <= to_signed(732,32);
				when 489 => sin_data_int <= to_signed(682,32); cos_data_int <= to_signed(731,32);
				when 490 => sin_data_int <= to_signed(683,32); cos_data_int <= to_signed(730,32);
				when 491 => sin_data_int <= to_signed(684,32); cos_data_int <= to_signed(728,32);
				when 492 => sin_data_int <= to_signed(685,32); cos_data_int <= to_signed(727,32);
				when 493 => sin_data_int <= to_signed(686,32); cos_data_int <= to_signed(726,32);
				when 494 => sin_data_int <= to_signed(687,32); cos_data_int <= to_signed(725,32);
				when 495 => sin_data_int <= to_signed(688,32); cos_data_int <= to_signed(724,32);
				when 496 => sin_data_int <= to_signed(690,32); cos_data_int <= to_signed(723,32);
				when 497 => sin_data_int <= to_signed(691,32); cos_data_int <= to_signed(722,32);
				when 498 => sin_data_int <= to_signed(692,32); cos_data_int <= to_signed(721,32);
				when 499 => sin_data_int <= to_signed(693,32); cos_data_int <= to_signed(720,32);
				when 500 => sin_data_int <= to_signed(694,32); cos_data_int <= to_signed(719,32);
				when 501 => sin_data_int <= to_signed(695,32); cos_data_int <= to_signed(718,32);
				when 502 => sin_data_int <= to_signed(696,32); cos_data_int <= to_signed(717,32);
				when 503 => sin_data_int <= to_signed(697,32); cos_data_int <= to_signed(716,32);
				when 504 => sin_data_int <= to_signed(698,32); cos_data_int <= to_signed(715,32);
				when 505 => sin_data_int <= to_signed(699,32); cos_data_int <= to_signed(714,32);
				when 506 => sin_data_int <= to_signed(701,32); cos_data_int <= to_signed(713,32);
				when 507 => sin_data_int <= to_signed(702,32); cos_data_int <= to_signed(711,32);
				when 508 => sin_data_int <= to_signed(703,32); cos_data_int <= to_signed(710,32);
				when 509 => sin_data_int <= to_signed(704,32); cos_data_int <= to_signed(709,32);
				when 510 => sin_data_int <= to_signed(705,32); cos_data_int <= to_signed(708,32);
				when 511 => sin_data_int <= to_signed(706,32); cos_data_int <= to_signed(707,32);
				when 512 => sin_data_int <= to_signed(707,32); cos_data_int <= to_signed(706,32);
				when 513 => sin_data_int <= to_signed(708,32); cos_data_int <= to_signed(705,32);
				when 514 => sin_data_int <= to_signed(709,32); cos_data_int <= to_signed(704,32);
				when 515 => sin_data_int <= to_signed(710,32); cos_data_int <= to_signed(703,32);
				when 516 => sin_data_int <= to_signed(711,32); cos_data_int <= to_signed(702,32);
				when 517 => sin_data_int <= to_signed(713,32); cos_data_int <= to_signed(701,32);
				when 518 => sin_data_int <= to_signed(714,32); cos_data_int <= to_signed(699,32);
				when 519 => sin_data_int <= to_signed(715,32); cos_data_int <= to_signed(698,32);
				when 520 => sin_data_int <= to_signed(716,32); cos_data_int <= to_signed(697,32);
				when 521 => sin_data_int <= to_signed(717,32); cos_data_int <= to_signed(696,32);
				when 522 => sin_data_int <= to_signed(718,32); cos_data_int <= to_signed(695,32);
				when 523 => sin_data_int <= to_signed(719,32); cos_data_int <= to_signed(694,32);
				when 524 => sin_data_int <= to_signed(720,32); cos_data_int <= to_signed(693,32);
				when 525 => sin_data_int <= to_signed(721,32); cos_data_int <= to_signed(692,32);
				when 526 => sin_data_int <= to_signed(722,32); cos_data_int <= to_signed(691,32);
				when 527 => sin_data_int <= to_signed(723,32); cos_data_int <= to_signed(690,32);
				when 528 => sin_data_int <= to_signed(724,32); cos_data_int <= to_signed(688,32);
				when 529 => sin_data_int <= to_signed(725,32); cos_data_int <= to_signed(687,32);
				when 530 => sin_data_int <= to_signed(726,32); cos_data_int <= to_signed(686,32);
				when 531 => sin_data_int <= to_signed(727,32); cos_data_int <= to_signed(685,32);
				when 532 => sin_data_int <= to_signed(728,32); cos_data_int <= to_signed(684,32);
				when 533 => sin_data_int <= to_signed(730,32); cos_data_int <= to_signed(683,32);
				when 534 => sin_data_int <= to_signed(731,32); cos_data_int <= to_signed(682,32);
				when 535 => sin_data_int <= to_signed(732,32); cos_data_int <= to_signed(681,32);
				when 536 => sin_data_int <= to_signed(733,32); cos_data_int <= to_signed(679,32);
				when 537 => sin_data_int <= to_signed(734,32); cos_data_int <= to_signed(678,32);
				when 538 => sin_data_int <= to_signed(735,32); cos_data_int <= to_signed(677,32);
				when 539 => sin_data_int <= to_signed(736,32); cos_data_int <= to_signed(676,32);
				when 540 => sin_data_int <= to_signed(737,32); cos_data_int <= to_signed(675,32);
				when 541 => sin_data_int <= to_signed(738,32); cos_data_int <= to_signed(674,32);
				when 542 => sin_data_int <= to_signed(739,32); cos_data_int <= to_signed(673,32);
				when 543 => sin_data_int <= to_signed(740,32); cos_data_int <= to_signed(672,32);
				when 544 => sin_data_int <= to_signed(741,32); cos_data_int <= to_signed(670,32);
				when 545 => sin_data_int <= to_signed(742,32); cos_data_int <= to_signed(669,32);
				when 546 => sin_data_int <= to_signed(743,32); cos_data_int <= to_signed(668,32);
				when 547 => sin_data_int <= to_signed(744,32); cos_data_int <= to_signed(667,32);
				when 548 => sin_data_int <= to_signed(745,32); cos_data_int <= to_signed(666,32);
				when 549 => sin_data_int <= to_signed(746,32); cos_data_int <= to_signed(665,32);
				when 550 => sin_data_int <= to_signed(747,32); cos_data_int <= to_signed(664,32);
				when 551 => sin_data_int <= to_signed(748,32); cos_data_int <= to_signed(662,32);
				when 552 => sin_data_int <= to_signed(749,32); cos_data_int <= to_signed(661,32);
				when 553 => sin_data_int <= to_signed(750,32); cos_data_int <= to_signed(660,32);
				when 554 => sin_data_int <= to_signed(751,32); cos_data_int <= to_signed(659,32);
				when 555 => sin_data_int <= to_signed(752,32); cos_data_int <= to_signed(658,32);
				when 556 => sin_data_int <= to_signed(753,32); cos_data_int <= to_signed(657,32);
				when 557 => sin_data_int <= to_signed(754,32); cos_data_int <= to_signed(655,32);
				when 558 => sin_data_int <= to_signed(755,32); cos_data_int <= to_signed(654,32);
				when 559 => sin_data_int <= to_signed(756,32); cos_data_int <= to_signed(653,32);
				when 560 => sin_data_int <= to_signed(757,32); cos_data_int <= to_signed(652,32);
				when 561 => sin_data_int <= to_signed(758,32); cos_data_int <= to_signed(651,32);
				when 562 => sin_data_int <= to_signed(759,32); cos_data_int <= to_signed(650,32);
				when 563 => sin_data_int <= to_signed(760,32); cos_data_int <= to_signed(649,32);
				when 564 => sin_data_int <= to_signed(761,32); cos_data_int <= to_signed(647,32);
				when 565 => sin_data_int <= to_signed(762,32); cos_data_int <= to_signed(646,32);
				when 566 => sin_data_int <= to_signed(763,32); cos_data_int <= to_signed(645,32);
				when 567 => sin_data_int <= to_signed(764,32); cos_data_int <= to_signed(644,32);
				when 568 => sin_data_int <= to_signed(765,32); cos_data_int <= to_signed(643,32);
				when 569 => sin_data_int <= to_signed(766,32); cos_data_int <= to_signed(641,32);
				when 570 => sin_data_int <= to_signed(767,32); cos_data_int <= to_signed(640,32);
				when 571 => sin_data_int <= to_signed(768,32); cos_data_int <= to_signed(639,32);
				when 572 => sin_data_int <= to_signed(769,32); cos_data_int <= to_signed(638,32);
				when 573 => sin_data_int <= to_signed(770,32); cos_data_int <= to_signed(637,32);
				when 574 => sin_data_int <= to_signed(771,32); cos_data_int <= to_signed(636,32);
				when 575 => sin_data_int <= to_signed(772,32); cos_data_int <= to_signed(634,32);
				when 576 => sin_data_int <= to_signed(773,32); cos_data_int <= to_signed(633,32);
				when 577 => sin_data_int <= to_signed(774,32); cos_data_int <= to_signed(632,32);
				when 578 => sin_data_int <= to_signed(775,32); cos_data_int <= to_signed(631,32);
				when 579 => sin_data_int <= to_signed(776,32); cos_data_int <= to_signed(630,32);
				when 580 => sin_data_int <= to_signed(777,32); cos_data_int <= to_signed(628,32);
				when 581 => sin_data_int <= to_signed(778,32); cos_data_int <= to_signed(627,32);
				when 582 => sin_data_int <= to_signed(779,32); cos_data_int <= to_signed(626,32);
				when 583 => sin_data_int <= to_signed(780,32); cos_data_int <= to_signed(625,32);
				when 584 => sin_data_int <= to_signed(781,32); cos_data_int <= to_signed(624,32);
				when 585 => sin_data_int <= to_signed(782,32); cos_data_int <= to_signed(622,32);
				when 586 => sin_data_int <= to_signed(783,32); cos_data_int <= to_signed(621,32);
				when 587 => sin_data_int <= to_signed(784,32); cos_data_int <= to_signed(620,32);
				when 588 => sin_data_int <= to_signed(785,32); cos_data_int <= to_signed(619,32);
				when 589 => sin_data_int <= to_signed(786,32); cos_data_int <= to_signed(618,32);
				when 590 => sin_data_int <= to_signed(786,32); cos_data_int <= to_signed(616,32);
				when 591 => sin_data_int <= to_signed(787,32); cos_data_int <= to_signed(615,32);
				when 592 => sin_data_int <= to_signed(788,32); cos_data_int <= to_signed(614,32);
				when 593 => sin_data_int <= to_signed(789,32); cos_data_int <= to_signed(613,32);
				when 594 => sin_data_int <= to_signed(790,32); cos_data_int <= to_signed(612,32);
				when 595 => sin_data_int <= to_signed(791,32); cos_data_int <= to_signed(610,32);
				when 596 => sin_data_int <= to_signed(792,32); cos_data_int <= to_signed(609,32);
				when 597 => sin_data_int <= to_signed(793,32); cos_data_int <= to_signed(608,32);
				when 598 => sin_data_int <= to_signed(794,32); cos_data_int <= to_signed(607,32);
				when 599 => sin_data_int <= to_signed(795,32); cos_data_int <= to_signed(606,32);
				when 600 => sin_data_int <= to_signed(796,32); cos_data_int <= to_signed(604,32);
				when 601 => sin_data_int <= to_signed(797,32); cos_data_int <= to_signed(603,32);
				when 602 => sin_data_int <= to_signed(798,32); cos_data_int <= to_signed(602,32);
				when 603 => sin_data_int <= to_signed(799,32); cos_data_int <= to_signed(601,32);
				when 604 => sin_data_int <= to_signed(800,32); cos_data_int <= to_signed(599,32);
				when 605 => sin_data_int <= to_signed(800,32); cos_data_int <= to_signed(598,32);
				when 606 => sin_data_int <= to_signed(801,32); cos_data_int <= to_signed(597,32);
				when 607 => sin_data_int <= to_signed(802,32); cos_data_int <= to_signed(596,32);
				when 608 => sin_data_int <= to_signed(803,32); cos_data_int <= to_signed(594,32);
				when 609 => sin_data_int <= to_signed(804,32); cos_data_int <= to_signed(593,32);
				when 610 => sin_data_int <= to_signed(805,32); cos_data_int <= to_signed(592,32);
				when 611 => sin_data_int <= to_signed(806,32); cos_data_int <= to_signed(591,32);
				when 612 => sin_data_int <= to_signed(807,32); cos_data_int <= to_signed(590,32);
				when 613 => sin_data_int <= to_signed(808,32); cos_data_int <= to_signed(588,32);
				when 614 => sin_data_int <= to_signed(809,32); cos_data_int <= to_signed(587,32);
				when 615 => sin_data_int <= to_signed(810,32); cos_data_int <= to_signed(586,32);
				when 616 => sin_data_int <= to_signed(810,32); cos_data_int <= to_signed(585,32);
				when 617 => sin_data_int <= to_signed(811,32); cos_data_int <= to_signed(583,32);
				when 618 => sin_data_int <= to_signed(812,32); cos_data_int <= to_signed(582,32);
				when 619 => sin_data_int <= to_signed(813,32); cos_data_int <= to_signed(581,32);
				when 620 => sin_data_int <= to_signed(814,32); cos_data_int <= to_signed(580,32);
				when 621 => sin_data_int <= to_signed(815,32); cos_data_int <= to_signed(578,32);
				when 622 => sin_data_int <= to_signed(816,32); cos_data_int <= to_signed(577,32);
				when 623 => sin_data_int <= to_signed(817,32); cos_data_int <= to_signed(576,32);
				when 624 => sin_data_int <= to_signed(818,32); cos_data_int <= to_signed(575,32);
				when 625 => sin_data_int <= to_signed(818,32); cos_data_int <= to_signed(573,32);
				when 626 => sin_data_int <= to_signed(819,32); cos_data_int <= to_signed(572,32);
				when 627 => sin_data_int <= to_signed(820,32); cos_data_int <= to_signed(571,32);
				when 628 => sin_data_int <= to_signed(821,32); cos_data_int <= to_signed(570,32);
				when 629 => sin_data_int <= to_signed(822,32); cos_data_int <= to_signed(568,32);
				when 630 => sin_data_int <= to_signed(823,32); cos_data_int <= to_signed(567,32);
				when 631 => sin_data_int <= to_signed(824,32); cos_data_int <= to_signed(566,32);
				when 632 => sin_data_int <= to_signed(825,32); cos_data_int <= to_signed(564,32);
				when 633 => sin_data_int <= to_signed(825,32); cos_data_int <= to_signed(563,32);
				when 634 => sin_data_int <= to_signed(826,32); cos_data_int <= to_signed(562,32);
				when 635 => sin_data_int <= to_signed(827,32); cos_data_int <= to_signed(561,32);
				when 636 => sin_data_int <= to_signed(828,32); cos_data_int <= to_signed(559,32);
				when 637 => sin_data_int <= to_signed(829,32); cos_data_int <= to_signed(558,32);
				when 638 => sin_data_int <= to_signed(830,32); cos_data_int <= to_signed(557,32);
				when 639 => sin_data_int <= to_signed(831,32); cos_data_int <= to_signed(556,32);
				when 640 => sin_data_int <= to_signed(831,32); cos_data_int <= to_signed(554,32);
				when 641 => sin_data_int <= to_signed(832,32); cos_data_int <= to_signed(553,32);
				when 642 => sin_data_int <= to_signed(833,32); cos_data_int <= to_signed(552,32);
				when 643 => sin_data_int <= to_signed(834,32); cos_data_int <= to_signed(550,32);
				when 644 => sin_data_int <= to_signed(835,32); cos_data_int <= to_signed(549,32);
				when 645 => sin_data_int <= to_signed(836,32); cos_data_int <= to_signed(548,32);
				when 646 => sin_data_int <= to_signed(837,32); cos_data_int <= to_signed(547,32);
				when 647 => sin_data_int <= to_signed(837,32); cos_data_int <= to_signed(545,32);
				when 648 => sin_data_int <= to_signed(838,32); cos_data_int <= to_signed(544,32);
				when 649 => sin_data_int <= to_signed(839,32); cos_data_int <= to_signed(543,32);
				when 650 => sin_data_int <= to_signed(840,32); cos_data_int <= to_signed(541,32);
				when 651 => sin_data_int <= to_signed(841,32); cos_data_int <= to_signed(540,32);
				when 652 => sin_data_int <= to_signed(842,32); cos_data_int <= to_signed(539,32);
				when 653 => sin_data_int <= to_signed(842,32); cos_data_int <= to_signed(538,32);
				when 654 => sin_data_int <= to_signed(843,32); cos_data_int <= to_signed(536,32);
				when 655 => sin_data_int <= to_signed(844,32); cos_data_int <= to_signed(535,32);
				when 656 => sin_data_int <= to_signed(845,32); cos_data_int <= to_signed(534,32);
				when 657 => sin_data_int <= to_signed(846,32); cos_data_int <= to_signed(532,32);
				when 658 => sin_data_int <= to_signed(846,32); cos_data_int <= to_signed(531,32);
				when 659 => sin_data_int <= to_signed(847,32); cos_data_int <= to_signed(530,32);
				when 660 => sin_data_int <= to_signed(848,32); cos_data_int <= to_signed(529,32);
				when 661 => sin_data_int <= to_signed(849,32); cos_data_int <= to_signed(527,32);
				when 662 => sin_data_int <= to_signed(850,32); cos_data_int <= to_signed(526,32);
				when 663 => sin_data_int <= to_signed(851,32); cos_data_int <= to_signed(525,32);
				when 664 => sin_data_int <= to_signed(851,32); cos_data_int <= to_signed(523,32);
				when 665 => sin_data_int <= to_signed(852,32); cos_data_int <= to_signed(522,32);
				when 666 => sin_data_int <= to_signed(853,32); cos_data_int <= to_signed(521,32);
				when 667 => sin_data_int <= to_signed(854,32); cos_data_int <= to_signed(519,32);
				when 668 => sin_data_int <= to_signed(855,32); cos_data_int <= to_signed(518,32);
				when 669 => sin_data_int <= to_signed(855,32); cos_data_int <= to_signed(517,32);
				when 670 => sin_data_int <= to_signed(856,32); cos_data_int <= to_signed(515,32);
				when 671 => sin_data_int <= to_signed(857,32); cos_data_int <= to_signed(514,32);
				when 672 => sin_data_int <= to_signed(858,32); cos_data_int <= to_signed(513,32);
				when 673 => sin_data_int <= to_signed(859,32); cos_data_int <= to_signed(511,32);
				when 674 => sin_data_int <= to_signed(859,32); cos_data_int <= to_signed(510,32);
				when 675 => sin_data_int <= to_signed(860,32); cos_data_int <= to_signed(509,32);
				when 676 => sin_data_int <= to_signed(861,32); cos_data_int <= to_signed(508,32);
				when 677 => sin_data_int <= to_signed(862,32); cos_data_int <= to_signed(506,32);
				when 678 => sin_data_int <= to_signed(862,32); cos_data_int <= to_signed(505,32);
				when 679 => sin_data_int <= to_signed(863,32); cos_data_int <= to_signed(504,32);
				when 680 => sin_data_int <= to_signed(864,32); cos_data_int <= to_signed(502,32);
				when 681 => sin_data_int <= to_signed(865,32); cos_data_int <= to_signed(501,32);
				when 682 => sin_data_int <= to_signed(866,32); cos_data_int <= to_signed(500,32);
				when 683 => sin_data_int <= to_signed(866,32); cos_data_int <= to_signed(498,32);
				when 684 => sin_data_int <= to_signed(867,32); cos_data_int <= to_signed(497,32);
				when 685 => sin_data_int <= to_signed(868,32); cos_data_int <= to_signed(496,32);
				when 686 => sin_data_int <= to_signed(869,32); cos_data_int <= to_signed(494,32);
				when 687 => sin_data_int <= to_signed(869,32); cos_data_int <= to_signed(493,32);
				when 688 => sin_data_int <= to_signed(870,32); cos_data_int <= to_signed(492,32);
				when 689 => sin_data_int <= to_signed(871,32); cos_data_int <= to_signed(490,32);
				when 690 => sin_data_int <= to_signed(872,32); cos_data_int <= to_signed(489,32);
				when 691 => sin_data_int <= to_signed(872,32); cos_data_int <= to_signed(488,32);
				when 692 => sin_data_int <= to_signed(873,32); cos_data_int <= to_signed(486,32);
				when 693 => sin_data_int <= to_signed(874,32); cos_data_int <= to_signed(485,32);
				when 694 => sin_data_int <= to_signed(875,32); cos_data_int <= to_signed(484,32);
				when 695 => sin_data_int <= to_signed(875,32); cos_data_int <= to_signed(482,32);
				when 696 => sin_data_int <= to_signed(876,32); cos_data_int <= to_signed(481,32);
				when 697 => sin_data_int <= to_signed(877,32); cos_data_int <= to_signed(479,32);
				when 698 => sin_data_int <= to_signed(878,32); cos_data_int <= to_signed(478,32);
				when 699 => sin_data_int <= to_signed(878,32); cos_data_int <= to_signed(477,32);
				when 700 => sin_data_int <= to_signed(879,32); cos_data_int <= to_signed(475,32);
				when 701 => sin_data_int <= to_signed(880,32); cos_data_int <= to_signed(474,32);
				when 702 => sin_data_int <= to_signed(880,32); cos_data_int <= to_signed(473,32);
				when 703 => sin_data_int <= to_signed(881,32); cos_data_int <= to_signed(471,32);
				when 704 => sin_data_int <= to_signed(882,32); cos_data_int <= to_signed(470,32);
				when 705 => sin_data_int <= to_signed(883,32); cos_data_int <= to_signed(469,32);
				when 706 => sin_data_int <= to_signed(883,32); cos_data_int <= to_signed(467,32);
				when 707 => sin_data_int <= to_signed(884,32); cos_data_int <= to_signed(466,32);
				when 708 => sin_data_int <= to_signed(885,32); cos_data_int <= to_signed(465,32);
				when 709 => sin_data_int <= to_signed(886,32); cos_data_int <= to_signed(463,32);
				when 710 => sin_data_int <= to_signed(886,32); cos_data_int <= to_signed(462,32);
				when 711 => sin_data_int <= to_signed(887,32); cos_data_int <= to_signed(461,32);
				when 712 => sin_data_int <= to_signed(888,32); cos_data_int <= to_signed(459,32);
				when 713 => sin_data_int <= to_signed(888,32); cos_data_int <= to_signed(458,32);
				when 714 => sin_data_int <= to_signed(889,32); cos_data_int <= to_signed(456,32);
				when 715 => sin_data_int <= to_signed(890,32); cos_data_int <= to_signed(455,32);
				when 716 => sin_data_int <= to_signed(890,32); cos_data_int <= to_signed(454,32);
				when 717 => sin_data_int <= to_signed(891,32); cos_data_int <= to_signed(452,32);
				when 718 => sin_data_int <= to_signed(892,32); cos_data_int <= to_signed(451,32);
				when 719 => sin_data_int <= to_signed(893,32); cos_data_int <= to_signed(450,32);
				when 720 => sin_data_int <= to_signed(893,32); cos_data_int <= to_signed(448,32);
				when 721 => sin_data_int <= to_signed(894,32); cos_data_int <= to_signed(447,32);
				when 722 => sin_data_int <= to_signed(895,32); cos_data_int <= to_signed(445,32);
				when 723 => sin_data_int <= to_signed(895,32); cos_data_int <= to_signed(444,32);
				when 724 => sin_data_int <= to_signed(896,32); cos_data_int <= to_signed(443,32);
				when 725 => sin_data_int <= to_signed(897,32); cos_data_int <= to_signed(441,32);
				when 726 => sin_data_int <= to_signed(897,32); cos_data_int <= to_signed(440,32);
				when 727 => sin_data_int <= to_signed(898,32); cos_data_int <= to_signed(439,32);
				when 728 => sin_data_int <= to_signed(899,32); cos_data_int <= to_signed(437,32);
				when 729 => sin_data_int <= to_signed(899,32); cos_data_int <= to_signed(436,32);
				when 730 => sin_data_int <= to_signed(900,32); cos_data_int <= to_signed(434,32);
				when 731 => sin_data_int <= to_signed(901,32); cos_data_int <= to_signed(433,32);
				when 732 => sin_data_int <= to_signed(901,32); cos_data_int <= to_signed(432,32);
				when 733 => sin_data_int <= to_signed(902,32); cos_data_int <= to_signed(430,32);
				when 734 => sin_data_int <= to_signed(903,32); cos_data_int <= to_signed(429,32);
				when 735 => sin_data_int <= to_signed(903,32); cos_data_int <= to_signed(428,32);
				when 736 => sin_data_int <= to_signed(904,32); cos_data_int <= to_signed(426,32);
				when 737 => sin_data_int <= to_signed(905,32); cos_data_int <= to_signed(425,32);
				when 738 => sin_data_int <= to_signed(905,32); cos_data_int <= to_signed(423,32);
				when 739 => sin_data_int <= to_signed(906,32); cos_data_int <= to_signed(422,32);
				when 740 => sin_data_int <= to_signed(907,32); cos_data_int <= to_signed(421,32);
				when 741 => sin_data_int <= to_signed(907,32); cos_data_int <= to_signed(419,32);
				when 742 => sin_data_int <= to_signed(908,32); cos_data_int <= to_signed(418,32);
				when 743 => sin_data_int <= to_signed(909,32); cos_data_int <= to_signed(416,32);
				when 744 => sin_data_int <= to_signed(909,32); cos_data_int <= to_signed(415,32);
				when 745 => sin_data_int <= to_signed(910,32); cos_data_int <= to_signed(414,32);
				when 746 => sin_data_int <= to_signed(910,32); cos_data_int <= to_signed(412,32);
				when 747 => sin_data_int <= to_signed(911,32); cos_data_int <= to_signed(411,32);
				when 748 => sin_data_int <= to_signed(912,32); cos_data_int <= to_signed(409,32);
				when 749 => sin_data_int <= to_signed(912,32); cos_data_int <= to_signed(408,32);
				when 750 => sin_data_int <= to_signed(913,32); cos_data_int <= to_signed(407,32);
				when 751 => sin_data_int <= to_signed(914,32); cos_data_int <= to_signed(405,32);
				when 752 => sin_data_int <= to_signed(914,32); cos_data_int <= to_signed(404,32);
				when 753 => sin_data_int <= to_signed(915,32); cos_data_int <= to_signed(402,32);
				when 754 => sin_data_int <= to_signed(915,32); cos_data_int <= to_signed(401,32);
				when 755 => sin_data_int <= to_signed(916,32); cos_data_int <= to_signed(400,32);
				when 756 => sin_data_int <= to_signed(917,32); cos_data_int <= to_signed(398,32);
				when 757 => sin_data_int <= to_signed(917,32); cos_data_int <= to_signed(397,32);
				when 758 => sin_data_int <= to_signed(918,32); cos_data_int <= to_signed(395,32);
				when 759 => sin_data_int <= to_signed(919,32); cos_data_int <= to_signed(394,32);
				when 760 => sin_data_int <= to_signed(919,32); cos_data_int <= to_signed(393,32);
				when 761 => sin_data_int <= to_signed(920,32); cos_data_int <= to_signed(391,32);
				when 762 => sin_data_int <= to_signed(920,32); cos_data_int <= to_signed(390,32);
				when 763 => sin_data_int <= to_signed(921,32); cos_data_int <= to_signed(388,32);
				when 764 => sin_data_int <= to_signed(922,32); cos_data_int <= to_signed(387,32);
				when 765 => sin_data_int <= to_signed(922,32); cos_data_int <= to_signed(386,32);
				when 766 => sin_data_int <= to_signed(923,32); cos_data_int <= to_signed(384,32);
				when 767 => sin_data_int <= to_signed(923,32); cos_data_int <= to_signed(383,32);
				when 768 => sin_data_int <= to_signed(924,32); cos_data_int <= to_signed(381,32);
				when 769 => sin_data_int <= to_signed(924,32); cos_data_int <= to_signed(380,32);
				when 770 => sin_data_int <= to_signed(925,32); cos_data_int <= to_signed(378,32);
				when 771 => sin_data_int <= to_signed(926,32); cos_data_int <= to_signed(377,32);
				when 772 => sin_data_int <= to_signed(926,32); cos_data_int <= to_signed(376,32);
				when 773 => sin_data_int <= to_signed(927,32); cos_data_int <= to_signed(374,32);
				when 774 => sin_data_int <= to_signed(927,32); cos_data_int <= to_signed(373,32);
				when 775 => sin_data_int <= to_signed(928,32); cos_data_int <= to_signed(371,32);
				when 776 => sin_data_int <= to_signed(929,32); cos_data_int <= to_signed(370,32);
				when 777 => sin_data_int <= to_signed(929,32); cos_data_int <= to_signed(368,32);
				when 778 => sin_data_int <= to_signed(930,32); cos_data_int <= to_signed(367,32);
				when 779 => sin_data_int <= to_signed(930,32); cos_data_int <= to_signed(366,32);
				when 780 => sin_data_int <= to_signed(931,32); cos_data_int <= to_signed(364,32);
				when 781 => sin_data_int <= to_signed(931,32); cos_data_int <= to_signed(363,32);
				when 782 => sin_data_int <= to_signed(932,32); cos_data_int <= to_signed(361,32);
				when 783 => sin_data_int <= to_signed(932,32); cos_data_int <= to_signed(360,32);
				when 784 => sin_data_int <= to_signed(933,32); cos_data_int <= to_signed(358,32);
				when 785 => sin_data_int <= to_signed(934,32); cos_data_int <= to_signed(357,32);
				when 786 => sin_data_int <= to_signed(934,32); cos_data_int <= to_signed(356,32);
				when 787 => sin_data_int <= to_signed(935,32); cos_data_int <= to_signed(354,32);
				when 788 => sin_data_int <= to_signed(935,32); cos_data_int <= to_signed(353,32);
				when 789 => sin_data_int <= to_signed(936,32); cos_data_int <= to_signed(351,32);
				when 790 => sin_data_int <= to_signed(936,32); cos_data_int <= to_signed(350,32);
				when 791 => sin_data_int <= to_signed(937,32); cos_data_int <= to_signed(348,32);
				when 792 => sin_data_int <= to_signed(937,32); cos_data_int <= to_signed(347,32);
				when 793 => sin_data_int <= to_signed(938,32); cos_data_int <= to_signed(346,32);
				when 794 => sin_data_int <= to_signed(938,32); cos_data_int <= to_signed(344,32);
				when 795 => sin_data_int <= to_signed(939,32); cos_data_int <= to_signed(343,32);
				when 796 => sin_data_int <= to_signed(939,32); cos_data_int <= to_signed(341,32);
				when 797 => sin_data_int <= to_signed(940,32); cos_data_int <= to_signed(340,32);
				when 798 => sin_data_int <= to_signed(941,32); cos_data_int <= to_signed(338,32);
				when 799 => sin_data_int <= to_signed(941,32); cos_data_int <= to_signed(337,32);
				when 800 => sin_data_int <= to_signed(942,32); cos_data_int <= to_signed(335,32);
				when 801 => sin_data_int <= to_signed(942,32); cos_data_int <= to_signed(334,32);
				when 802 => sin_data_int <= to_signed(943,32); cos_data_int <= to_signed(333,32);
				when 803 => sin_data_int <= to_signed(943,32); cos_data_int <= to_signed(331,32);
				when 804 => sin_data_int <= to_signed(944,32); cos_data_int <= to_signed(330,32);
				when 805 => sin_data_int <= to_signed(944,32); cos_data_int <= to_signed(328,32);
				when 806 => sin_data_int <= to_signed(945,32); cos_data_int <= to_signed(327,32);
				when 807 => sin_data_int <= to_signed(945,32); cos_data_int <= to_signed(325,32);
				when 808 => sin_data_int <= to_signed(946,32); cos_data_int <= to_signed(324,32);
				when 809 => sin_data_int <= to_signed(946,32); cos_data_int <= to_signed(322,32);
				when 810 => sin_data_int <= to_signed(947,32); cos_data_int <= to_signed(321,32);
				when 811 => sin_data_int <= to_signed(947,32); cos_data_int <= to_signed(320,32);
				when 812 => sin_data_int <= to_signed(948,32); cos_data_int <= to_signed(318,32);
				when 813 => sin_data_int <= to_signed(948,32); cos_data_int <= to_signed(317,32);
				when 814 => sin_data_int <= to_signed(949,32); cos_data_int <= to_signed(315,32);
				when 815 => sin_data_int <= to_signed(949,32); cos_data_int <= to_signed(314,32);
				when 816 => sin_data_int <= to_signed(950,32); cos_data_int <= to_signed(312,32);
				when 817 => sin_data_int <= to_signed(950,32); cos_data_int <= to_signed(311,32);
				when 818 => sin_data_int <= to_signed(950,32); cos_data_int <= to_signed(309,32);
				when 819 => sin_data_int <= to_signed(951,32); cos_data_int <= to_signed(308,32);
				when 820 => sin_data_int <= to_signed(951,32); cos_data_int <= to_signed(306,32);
				when 821 => sin_data_int <= to_signed(952,32); cos_data_int <= to_signed(305,32);
				when 822 => sin_data_int <= to_signed(952,32); cos_data_int <= to_signed(303,32);
				when 823 => sin_data_int <= to_signed(953,32); cos_data_int <= to_signed(302,32);
				when 824 => sin_data_int <= to_signed(953,32); cos_data_int <= to_signed(301,32);
				when 825 => sin_data_int <= to_signed(954,32); cos_data_int <= to_signed(299,32);
				when 826 => sin_data_int <= to_signed(954,32); cos_data_int <= to_signed(298,32);
				when 827 => sin_data_int <= to_signed(955,32); cos_data_int <= to_signed(296,32);
				when 828 => sin_data_int <= to_signed(955,32); cos_data_int <= to_signed(295,32);
				when 829 => sin_data_int <= to_signed(956,32); cos_data_int <= to_signed(293,32);
				when 830 => sin_data_int <= to_signed(956,32); cos_data_int <= to_signed(292,32);
				when 831 => sin_data_int <= to_signed(956,32); cos_data_int <= to_signed(290,32);
				when 832 => sin_data_int <= to_signed(957,32); cos_data_int <= to_signed(289,32);
				when 833 => sin_data_int <= to_signed(957,32); cos_data_int <= to_signed(287,32);
				when 834 => sin_data_int <= to_signed(958,32); cos_data_int <= to_signed(286,32);
				when 835 => sin_data_int <= to_signed(958,32); cos_data_int <= to_signed(284,32);
				when 836 => sin_data_int <= to_signed(959,32); cos_data_int <= to_signed(283,32);
				when 837 => sin_data_int <= to_signed(959,32); cos_data_int <= to_signed(281,32);
				when 838 => sin_data_int <= to_signed(960,32); cos_data_int <= to_signed(280,32);
				when 839 => sin_data_int <= to_signed(960,32); cos_data_int <= to_signed(279,32);
				when 840 => sin_data_int <= to_signed(960,32); cos_data_int <= to_signed(277,32);
				when 841 => sin_data_int <= to_signed(961,32); cos_data_int <= to_signed(276,32);
				when 842 => sin_data_int <= to_signed(961,32); cos_data_int <= to_signed(274,32);
				when 843 => sin_data_int <= to_signed(962,32); cos_data_int <= to_signed(273,32);
				when 844 => sin_data_int <= to_signed(962,32); cos_data_int <= to_signed(271,32);
				when 845 => sin_data_int <= to_signed(963,32); cos_data_int <= to_signed(270,32);
				when 846 => sin_data_int <= to_signed(963,32); cos_data_int <= to_signed(268,32);
				when 847 => sin_data_int <= to_signed(963,32); cos_data_int <= to_signed(267,32);
				when 848 => sin_data_int <= to_signed(964,32); cos_data_int <= to_signed(265,32);
				when 849 => sin_data_int <= to_signed(964,32); cos_data_int <= to_signed(264,32);
				when 850 => sin_data_int <= to_signed(965,32); cos_data_int <= to_signed(262,32);
				when 851 => sin_data_int <= to_signed(965,32); cos_data_int <= to_signed(261,32);
				when 852 => sin_data_int <= to_signed(965,32); cos_data_int <= to_signed(259,32);
				when 853 => sin_data_int <= to_signed(966,32); cos_data_int <= to_signed(258,32);
				when 854 => sin_data_int <= to_signed(966,32); cos_data_int <= to_signed(256,32);
				when 855 => sin_data_int <= to_signed(967,32); cos_data_int <= to_signed(255,32);
				when 856 => sin_data_int <= to_signed(967,32); cos_data_int <= to_signed(253,32);
				when 857 => sin_data_int <= to_signed(967,32); cos_data_int <= to_signed(252,32);
				when 858 => sin_data_int <= to_signed(968,32); cos_data_int <= to_signed(250,32);
				when 859 => sin_data_int <= to_signed(968,32); cos_data_int <= to_signed(249,32);
				when 860 => sin_data_int <= to_signed(969,32); cos_data_int <= to_signed(247,32);
				when 861 => sin_data_int <= to_signed(969,32); cos_data_int <= to_signed(246,32);
				when 862 => sin_data_int <= to_signed(969,32); cos_data_int <= to_signed(244,32);
				when 863 => sin_data_int <= to_signed(970,32); cos_data_int <= to_signed(243,32);
				when 864 => sin_data_int <= to_signed(970,32); cos_data_int <= to_signed(241,32);
				when 865 => sin_data_int <= to_signed(970,32); cos_data_int <= to_signed(240,32);
				when 866 => sin_data_int <= to_signed(971,32); cos_data_int <= to_signed(239,32);
				when 867 => sin_data_int <= to_signed(971,32); cos_data_int <= to_signed(237,32);
				when 868 => sin_data_int <= to_signed(972,32); cos_data_int <= to_signed(236,32);
				when 869 => sin_data_int <= to_signed(972,32); cos_data_int <= to_signed(234,32);
				when 870 => sin_data_int <= to_signed(972,32); cos_data_int <= to_signed(233,32);
				when 871 => sin_data_int <= to_signed(973,32); cos_data_int <= to_signed(231,32);
				when 872 => sin_data_int <= to_signed(973,32); cos_data_int <= to_signed(230,32);
				when 873 => sin_data_int <= to_signed(973,32); cos_data_int <= to_signed(228,32);
				when 874 => sin_data_int <= to_signed(974,32); cos_data_int <= to_signed(227,32);
				when 875 => sin_data_int <= to_signed(974,32); cos_data_int <= to_signed(225,32);
				when 876 => sin_data_int <= to_signed(974,32); cos_data_int <= to_signed(224,32);
				when 877 => sin_data_int <= to_signed(975,32); cos_data_int <= to_signed(222,32);
				when 878 => sin_data_int <= to_signed(975,32); cos_data_int <= to_signed(221,32);
				when 879 => sin_data_int <= to_signed(975,32); cos_data_int <= to_signed(219,32);
				when 880 => sin_data_int <= to_signed(976,32); cos_data_int <= to_signed(218,32);
				when 881 => sin_data_int <= to_signed(976,32); cos_data_int <= to_signed(216,32);
				when 882 => sin_data_int <= to_signed(976,32); cos_data_int <= to_signed(215,32);
				when 883 => sin_data_int <= to_signed(977,32); cos_data_int <= to_signed(213,32);
				when 884 => sin_data_int <= to_signed(977,32); cos_data_int <= to_signed(212,32);
				when 885 => sin_data_int <= to_signed(977,32); cos_data_int <= to_signed(210,32);
				when 886 => sin_data_int <= to_signed(978,32); cos_data_int <= to_signed(209,32);
				when 887 => sin_data_int <= to_signed(978,32); cos_data_int <= to_signed(207,32);
				when 888 => sin_data_int <= to_signed(978,32); cos_data_int <= to_signed(206,32);
				when 889 => sin_data_int <= to_signed(979,32); cos_data_int <= to_signed(204,32);
				when 890 => sin_data_int <= to_signed(979,32); cos_data_int <= to_signed(203,32);
				when 891 => sin_data_int <= to_signed(979,32); cos_data_int <= to_signed(201,32);
				when 892 => sin_data_int <= to_signed(980,32); cos_data_int <= to_signed(200,32);
				when 893 => sin_data_int <= to_signed(980,32); cos_data_int <= to_signed(198,32);
				when 894 => sin_data_int <= to_signed(980,32); cos_data_int <= to_signed(197,32);
				when 895 => sin_data_int <= to_signed(980,32); cos_data_int <= to_signed(195,32);
				when 896 => sin_data_int <= to_signed(981,32); cos_data_int <= to_signed(194,32);
				when 897 => sin_data_int <= to_signed(981,32); cos_data_int <= to_signed(192,32);
				when 898 => sin_data_int <= to_signed(981,32); cos_data_int <= to_signed(191,32);
				when 899 => sin_data_int <= to_signed(982,32); cos_data_int <= to_signed(189,32);
				when 900 => sin_data_int <= to_signed(982,32); cos_data_int <= to_signed(188,32);
				when 901 => sin_data_int <= to_signed(982,32); cos_data_int <= to_signed(186,32);
				when 902 => sin_data_int <= to_signed(983,32); cos_data_int <= to_signed(185,32);
				when 903 => sin_data_int <= to_signed(983,32); cos_data_int <= to_signed(183,32);
				when 904 => sin_data_int <= to_signed(983,32); cos_data_int <= to_signed(182,32);
				when 905 => sin_data_int <= to_signed(983,32); cos_data_int <= to_signed(180,32);
				when 906 => sin_data_int <= to_signed(984,32); cos_data_int <= to_signed(179,32);
				when 907 => sin_data_int <= to_signed(984,32); cos_data_int <= to_signed(177,32);
				when 908 => sin_data_int <= to_signed(984,32); cos_data_int <= to_signed(175,32);
				when 909 => sin_data_int <= to_signed(984,32); cos_data_int <= to_signed(174,32);
				when 910 => sin_data_int <= to_signed(985,32); cos_data_int <= to_signed(172,32);
				when 911 => sin_data_int <= to_signed(985,32); cos_data_int <= to_signed(171,32);
				when 912 => sin_data_int <= to_signed(985,32); cos_data_int <= to_signed(169,32);
				when 913 => sin_data_int <= to_signed(986,32); cos_data_int <= to_signed(168,32);
				when 914 => sin_data_int <= to_signed(986,32); cos_data_int <= to_signed(166,32);
				when 915 => sin_data_int <= to_signed(986,32); cos_data_int <= to_signed(165,32);
				when 916 => sin_data_int <= to_signed(986,32); cos_data_int <= to_signed(163,32);
				when 917 => sin_data_int <= to_signed(987,32); cos_data_int <= to_signed(162,32);
				when 918 => sin_data_int <= to_signed(987,32); cos_data_int <= to_signed(160,32);
				when 919 => sin_data_int <= to_signed(987,32); cos_data_int <= to_signed(159,32);
				when 920 => sin_data_int <= to_signed(987,32); cos_data_int <= to_signed(157,32);
				when 921 => sin_data_int <= to_signed(988,32); cos_data_int <= to_signed(156,32);
				when 922 => sin_data_int <= to_signed(988,32); cos_data_int <= to_signed(154,32);
				when 923 => sin_data_int <= to_signed(988,32); cos_data_int <= to_signed(153,32);
				when 924 => sin_data_int <= to_signed(988,32); cos_data_int <= to_signed(151,32);
				when 925 => sin_data_int <= to_signed(988,32); cos_data_int <= to_signed(150,32);
				when 926 => sin_data_int <= to_signed(989,32); cos_data_int <= to_signed(148,32);
				when 927 => sin_data_int <= to_signed(989,32); cos_data_int <= to_signed(147,32);
				when 928 => sin_data_int <= to_signed(989,32); cos_data_int <= to_signed(145,32);
				when 929 => sin_data_int <= to_signed(989,32); cos_data_int <= to_signed(144,32);
				when 930 => sin_data_int <= to_signed(990,32); cos_data_int <= to_signed(142,32);
				when 931 => sin_data_int <= to_signed(990,32); cos_data_int <= to_signed(141,32);
				when 932 => sin_data_int <= to_signed(990,32); cos_data_int <= to_signed(139,32);
				when 933 => sin_data_int <= to_signed(990,32); cos_data_int <= to_signed(138,32);
				when 934 => sin_data_int <= to_signed(990,32); cos_data_int <= to_signed(136,32);
				when 935 => sin_data_int <= to_signed(991,32); cos_data_int <= to_signed(135,32);
				when 936 => sin_data_int <= to_signed(991,32); cos_data_int <= to_signed(133,32);
				when 937 => sin_data_int <= to_signed(991,32); cos_data_int <= to_signed(132,32);
				when 938 => sin_data_int <= to_signed(991,32); cos_data_int <= to_signed(130,32);
				when 939 => sin_data_int <= to_signed(992,32); cos_data_int <= to_signed(128,32);
				when 940 => sin_data_int <= to_signed(992,32); cos_data_int <= to_signed(127,32);
				when 941 => sin_data_int <= to_signed(992,32); cos_data_int <= to_signed(125,32);
				when 942 => sin_data_int <= to_signed(992,32); cos_data_int <= to_signed(124,32);
				when 943 => sin_data_int <= to_signed(992,32); cos_data_int <= to_signed(122,32);
				when 944 => sin_data_int <= to_signed(992,32); cos_data_int <= to_signed(121,32);
				when 945 => sin_data_int <= to_signed(993,32); cos_data_int <= to_signed(119,32);
				when 946 => sin_data_int <= to_signed(993,32); cos_data_int <= to_signed(118,32);
				when 947 => sin_data_int <= to_signed(993,32); cos_data_int <= to_signed(116,32);
				when 948 => sin_data_int <= to_signed(993,32); cos_data_int <= to_signed(115,32);
				when 949 => sin_data_int <= to_signed(993,32); cos_data_int <= to_signed(113,32);
				when 950 => sin_data_int <= to_signed(994,32); cos_data_int <= to_signed(112,32);
				when 951 => sin_data_int <= to_signed(994,32); cos_data_int <= to_signed(110,32);
				when 952 => sin_data_int <= to_signed(994,32); cos_data_int <= to_signed(109,32);
				when 953 => sin_data_int <= to_signed(994,32); cos_data_int <= to_signed(107,32);
				when 954 => sin_data_int <= to_signed(994,32); cos_data_int <= to_signed(106,32);
				when 955 => sin_data_int <= to_signed(994,32); cos_data_int <= to_signed(104,32);
				when 956 => sin_data_int <= to_signed(995,32); cos_data_int <= to_signed(103,32);
				when 957 => sin_data_int <= to_signed(995,32); cos_data_int <= to_signed(101,32);
				when 958 => sin_data_int <= to_signed(995,32); cos_data_int <= to_signed(100,32);
				when 959 => sin_data_int <= to_signed(995,32); cos_data_int <= to_signed(98,32);
				when 960 => sin_data_int <= to_signed(995,32); cos_data_int <= to_signed(96,32);
				when 961 => sin_data_int <= to_signed(995,32); cos_data_int <= to_signed(95,32);
				when 962 => sin_data_int <= to_signed(995,32); cos_data_int <= to_signed(93,32);
				when 963 => sin_data_int <= to_signed(996,32); cos_data_int <= to_signed(92,32);
				when 964 => sin_data_int <= to_signed(996,32); cos_data_int <= to_signed(90,32);
				when 965 => sin_data_int <= to_signed(996,32); cos_data_int <= to_signed(89,32);
				when 966 => sin_data_int <= to_signed(996,32); cos_data_int <= to_signed(87,32);
				when 967 => sin_data_int <= to_signed(996,32); cos_data_int <= to_signed(86,32);
				when 968 => sin_data_int <= to_signed(996,32); cos_data_int <= to_signed(84,32);
				when 969 => sin_data_int <= to_signed(996,32); cos_data_int <= to_signed(83,32);
				when 970 => sin_data_int <= to_signed(997,32); cos_data_int <= to_signed(81,32);
				when 971 => sin_data_int <= to_signed(997,32); cos_data_int <= to_signed(80,32);
				when 972 => sin_data_int <= to_signed(997,32); cos_data_int <= to_signed(78,32);
				when 973 => sin_data_int <= to_signed(997,32); cos_data_int <= to_signed(77,32);
				when 974 => sin_data_int <= to_signed(997,32); cos_data_int <= to_signed(75,32);
				when 975 => sin_data_int <= to_signed(997,32); cos_data_int <= to_signed(74,32);
				when 976 => sin_data_int <= to_signed(997,32); cos_data_int <= to_signed(72,32);
				when 977 => sin_data_int <= to_signed(997,32); cos_data_int <= to_signed(71,32);
				when 978 => sin_data_int <= to_signed(998,32); cos_data_int <= to_signed(69,32);
				when 979 => sin_data_int <= to_signed(998,32); cos_data_int <= to_signed(67,32);
				when 980 => sin_data_int <= to_signed(998,32); cos_data_int <= to_signed(66,32);
				when 981 => sin_data_int <= to_signed(998,32); cos_data_int <= to_signed(64,32);
				when 982 => sin_data_int <= to_signed(998,32); cos_data_int <= to_signed(63,32);
				when 983 => sin_data_int <= to_signed(998,32); cos_data_int <= to_signed(61,32);
				when 984 => sin_data_int <= to_signed(998,32); cos_data_int <= to_signed(60,32);
				when 985 => sin_data_int <= to_signed(998,32); cos_data_int <= to_signed(58,32);
				when 986 => sin_data_int <= to_signed(998,32); cos_data_int <= to_signed(57,32);
				when 987 => sin_data_int <= to_signed(998,32); cos_data_int <= to_signed(55,32);
				when 988 => sin_data_int <= to_signed(998,32); cos_data_int <= to_signed(54,32);
				when 989 => sin_data_int <= to_signed(999,32); cos_data_int <= to_signed(52,32);
				when 990 => sin_data_int <= to_signed(999,32); cos_data_int <= to_signed(51,32);
				when 991 => sin_data_int <= to_signed(999,32); cos_data_int <= to_signed(49,32);
				when 992 => sin_data_int <= to_signed(999,32); cos_data_int <= to_signed(48,32);
				when 993 => sin_data_int <= to_signed(999,32); cos_data_int <= to_signed(46,32);
				when 994 => sin_data_int <= to_signed(999,32); cos_data_int <= to_signed(44,32);
				when 995 => sin_data_int <= to_signed(999,32); cos_data_int <= to_signed(43,32);
				when 996 => sin_data_int <= to_signed(999,32); cos_data_int <= to_signed(41,32);
				when 997 => sin_data_int <= to_signed(999,32); cos_data_int <= to_signed(40,32);
				when 998 => sin_data_int <= to_signed(999,32); cos_data_int <= to_signed(38,32);
				when 999 => sin_data_int <= to_signed(999,32); cos_data_int <= to_signed(37,32);
				when 1000 => sin_data_int <= to_signed(999,32); cos_data_int <= to_signed(35,32);
				when 1001 => sin_data_int <= to_signed(999,32); cos_data_int <= to_signed(34,32);
				when 1002 => sin_data_int <= to_signed(999,32); cos_data_int <= to_signed(32,32);
				when 1003 => sin_data_int <= to_signed(999,32); cos_data_int <= to_signed(31,32);
				when 1004 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(29,32);
				when 1005 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(28,32);
				when 1006 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(26,32);
				when 1007 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(25,32);
				when 1008 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(23,32);
				when 1009 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(21,32);
				when 1010 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(20,32);
				when 1011 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(18,32);
				when 1012 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(17,32);
				when 1013 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(15,32);
				when 1014 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(14,32);
				when 1015 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(12,32);
				when 1016 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(11,32);
				when 1017 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(9,32);
				when 1018 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(8,32);
				when 1019 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(6,32);
				when 1020 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(5,32);
				when 1021 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(3,32);
				when 1022 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(2,32);
				when 1023 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(0,32);
				when 1024 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(-2,32);
				when 1025 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(-3,32);
				when 1026 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(-5,32);
				when 1027 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(-6,32);
				when 1028 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(-8,32);
				when 1029 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(-9,32);
				when 1030 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(-11,32);
				when 1031 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(-12,32);
				when 1032 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(-14,32);
				when 1033 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(-15,32);
				when 1034 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(-17,32);
				when 1035 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(-18,32);
				when 1036 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(-20,32);
				when 1037 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(-21,32);
				when 1038 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(-23,32);
				when 1039 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(-25,32);
				when 1040 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(-26,32);
				when 1041 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(-28,32);
				when 1042 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(-29,32);
				when 1043 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(-31,32);
				when 1044 => sin_data_int <= to_signed(1000,32); cos_data_int <= to_signed(-32,32);
				when 1045 => sin_data_int <= to_signed(999,32); cos_data_int <= to_signed(-34,32);
				when 1046 => sin_data_int <= to_signed(999,32); cos_data_int <= to_signed(-35,32);
				when 1047 => sin_data_int <= to_signed(999,32); cos_data_int <= to_signed(-37,32);
				when 1048 => sin_data_int <= to_signed(999,32); cos_data_int <= to_signed(-38,32);
				when 1049 => sin_data_int <= to_signed(999,32); cos_data_int <= to_signed(-40,32);
				when 1050 => sin_data_int <= to_signed(999,32); cos_data_int <= to_signed(-41,32);
				when 1051 => sin_data_int <= to_signed(999,32); cos_data_int <= to_signed(-43,32);
				when 1052 => sin_data_int <= to_signed(999,32); cos_data_int <= to_signed(-44,32);
				when 1053 => sin_data_int <= to_signed(999,32); cos_data_int <= to_signed(-46,32);
				when 1054 => sin_data_int <= to_signed(999,32); cos_data_int <= to_signed(-48,32);
				when 1055 => sin_data_int <= to_signed(999,32); cos_data_int <= to_signed(-49,32);
				when 1056 => sin_data_int <= to_signed(999,32); cos_data_int <= to_signed(-51,32);
				when 1057 => sin_data_int <= to_signed(999,32); cos_data_int <= to_signed(-52,32);
				when 1058 => sin_data_int <= to_signed(999,32); cos_data_int <= to_signed(-54,32);
				when 1059 => sin_data_int <= to_signed(999,32); cos_data_int <= to_signed(-55,32);
				when 1060 => sin_data_int <= to_signed(998,32); cos_data_int <= to_signed(-57,32);
				when 1061 => sin_data_int <= to_signed(998,32); cos_data_int <= to_signed(-58,32);
				when 1062 => sin_data_int <= to_signed(998,32); cos_data_int <= to_signed(-60,32);
				when 1063 => sin_data_int <= to_signed(998,32); cos_data_int <= to_signed(-61,32);
				when 1064 => sin_data_int <= to_signed(998,32); cos_data_int <= to_signed(-63,32);
				when 1065 => sin_data_int <= to_signed(998,32); cos_data_int <= to_signed(-64,32);
				when 1066 => sin_data_int <= to_signed(998,32); cos_data_int <= to_signed(-66,32);
				when 1067 => sin_data_int <= to_signed(998,32); cos_data_int <= to_signed(-67,32);
				when 1068 => sin_data_int <= to_signed(998,32); cos_data_int <= to_signed(-69,32);
				when 1069 => sin_data_int <= to_signed(998,32); cos_data_int <= to_signed(-71,32);
				when 1070 => sin_data_int <= to_signed(998,32); cos_data_int <= to_signed(-72,32);
				when 1071 => sin_data_int <= to_signed(997,32); cos_data_int <= to_signed(-74,32);
				when 1072 => sin_data_int <= to_signed(997,32); cos_data_int <= to_signed(-75,32);
				when 1073 => sin_data_int <= to_signed(997,32); cos_data_int <= to_signed(-77,32);
				when 1074 => sin_data_int <= to_signed(997,32); cos_data_int <= to_signed(-78,32);
				when 1075 => sin_data_int <= to_signed(997,32); cos_data_int <= to_signed(-80,32);
				when 1076 => sin_data_int <= to_signed(997,32); cos_data_int <= to_signed(-81,32);
				when 1077 => sin_data_int <= to_signed(997,32); cos_data_int <= to_signed(-83,32);
				when 1078 => sin_data_int <= to_signed(997,32); cos_data_int <= to_signed(-84,32);
				when 1079 => sin_data_int <= to_signed(996,32); cos_data_int <= to_signed(-86,32);
				when 1080 => sin_data_int <= to_signed(996,32); cos_data_int <= to_signed(-87,32);
				when 1081 => sin_data_int <= to_signed(996,32); cos_data_int <= to_signed(-89,32);
				when 1082 => sin_data_int <= to_signed(996,32); cos_data_int <= to_signed(-90,32);
				when 1083 => sin_data_int <= to_signed(996,32); cos_data_int <= to_signed(-92,32);
				when 1084 => sin_data_int <= to_signed(996,32); cos_data_int <= to_signed(-93,32);
				when 1085 => sin_data_int <= to_signed(996,32); cos_data_int <= to_signed(-95,32);
				when 1086 => sin_data_int <= to_signed(995,32); cos_data_int <= to_signed(-96,32);
				when 1087 => sin_data_int <= to_signed(995,32); cos_data_int <= to_signed(-98,32);
				when 1088 => sin_data_int <= to_signed(995,32); cos_data_int <= to_signed(-100,32);
				when 1089 => sin_data_int <= to_signed(995,32); cos_data_int <= to_signed(-101,32);
				when 1090 => sin_data_int <= to_signed(995,32); cos_data_int <= to_signed(-103,32);
				when 1091 => sin_data_int <= to_signed(995,32); cos_data_int <= to_signed(-104,32);
				when 1092 => sin_data_int <= to_signed(995,32); cos_data_int <= to_signed(-106,32);
				when 1093 => sin_data_int <= to_signed(994,32); cos_data_int <= to_signed(-107,32);
				when 1094 => sin_data_int <= to_signed(994,32); cos_data_int <= to_signed(-109,32);
				when 1095 => sin_data_int <= to_signed(994,32); cos_data_int <= to_signed(-110,32);
				when 1096 => sin_data_int <= to_signed(994,32); cos_data_int <= to_signed(-112,32);
				when 1097 => sin_data_int <= to_signed(994,32); cos_data_int <= to_signed(-113,32);
				when 1098 => sin_data_int <= to_signed(994,32); cos_data_int <= to_signed(-115,32);
				when 1099 => sin_data_int <= to_signed(993,32); cos_data_int <= to_signed(-116,32);
				when 1100 => sin_data_int <= to_signed(993,32); cos_data_int <= to_signed(-118,32);
				when 1101 => sin_data_int <= to_signed(993,32); cos_data_int <= to_signed(-119,32);
				when 1102 => sin_data_int <= to_signed(993,32); cos_data_int <= to_signed(-121,32);
				when 1103 => sin_data_int <= to_signed(993,32); cos_data_int <= to_signed(-122,32);
				when 1104 => sin_data_int <= to_signed(992,32); cos_data_int <= to_signed(-124,32);
				when 1105 => sin_data_int <= to_signed(992,32); cos_data_int <= to_signed(-125,32);
				when 1106 => sin_data_int <= to_signed(992,32); cos_data_int <= to_signed(-127,32);
				when 1107 => sin_data_int <= to_signed(992,32); cos_data_int <= to_signed(-128,32);
				when 1108 => sin_data_int <= to_signed(992,32); cos_data_int <= to_signed(-130,32);
				when 1109 => sin_data_int <= to_signed(992,32); cos_data_int <= to_signed(-132,32);
				when 1110 => sin_data_int <= to_signed(991,32); cos_data_int <= to_signed(-133,32);
				when 1111 => sin_data_int <= to_signed(991,32); cos_data_int <= to_signed(-135,32);
				when 1112 => sin_data_int <= to_signed(991,32); cos_data_int <= to_signed(-136,32);
				when 1113 => sin_data_int <= to_signed(991,32); cos_data_int <= to_signed(-138,32);
				when 1114 => sin_data_int <= to_signed(990,32); cos_data_int <= to_signed(-139,32);
				when 1115 => sin_data_int <= to_signed(990,32); cos_data_int <= to_signed(-141,32);
				when 1116 => sin_data_int <= to_signed(990,32); cos_data_int <= to_signed(-142,32);
				when 1117 => sin_data_int <= to_signed(990,32); cos_data_int <= to_signed(-144,32);
				when 1118 => sin_data_int <= to_signed(990,32); cos_data_int <= to_signed(-145,32);
				when 1119 => sin_data_int <= to_signed(989,32); cos_data_int <= to_signed(-147,32);
				when 1120 => sin_data_int <= to_signed(989,32); cos_data_int <= to_signed(-148,32);
				when 1121 => sin_data_int <= to_signed(989,32); cos_data_int <= to_signed(-150,32);
				when 1122 => sin_data_int <= to_signed(989,32); cos_data_int <= to_signed(-151,32);
				when 1123 => sin_data_int <= to_signed(988,32); cos_data_int <= to_signed(-153,32);
				when 1124 => sin_data_int <= to_signed(988,32); cos_data_int <= to_signed(-154,32);
				when 1125 => sin_data_int <= to_signed(988,32); cos_data_int <= to_signed(-156,32);
				when 1126 => sin_data_int <= to_signed(988,32); cos_data_int <= to_signed(-157,32);
				when 1127 => sin_data_int <= to_signed(988,32); cos_data_int <= to_signed(-159,32);
				when 1128 => sin_data_int <= to_signed(987,32); cos_data_int <= to_signed(-160,32);
				when 1129 => sin_data_int <= to_signed(987,32); cos_data_int <= to_signed(-162,32);
				when 1130 => sin_data_int <= to_signed(987,32); cos_data_int <= to_signed(-163,32);
				when 1131 => sin_data_int <= to_signed(987,32); cos_data_int <= to_signed(-165,32);
				when 1132 => sin_data_int <= to_signed(986,32); cos_data_int <= to_signed(-166,32);
				when 1133 => sin_data_int <= to_signed(986,32); cos_data_int <= to_signed(-168,32);
				when 1134 => sin_data_int <= to_signed(986,32); cos_data_int <= to_signed(-169,32);
				when 1135 => sin_data_int <= to_signed(986,32); cos_data_int <= to_signed(-171,32);
				when 1136 => sin_data_int <= to_signed(985,32); cos_data_int <= to_signed(-172,32);
				when 1137 => sin_data_int <= to_signed(985,32); cos_data_int <= to_signed(-174,32);
				when 1138 => sin_data_int <= to_signed(985,32); cos_data_int <= to_signed(-175,32);
				when 1139 => sin_data_int <= to_signed(984,32); cos_data_int <= to_signed(-177,32);
				when 1140 => sin_data_int <= to_signed(984,32); cos_data_int <= to_signed(-179,32);
				when 1141 => sin_data_int <= to_signed(984,32); cos_data_int <= to_signed(-180,32);
				when 1142 => sin_data_int <= to_signed(984,32); cos_data_int <= to_signed(-182,32);
				when 1143 => sin_data_int <= to_signed(983,32); cos_data_int <= to_signed(-183,32);
				when 1144 => sin_data_int <= to_signed(983,32); cos_data_int <= to_signed(-185,32);
				when 1145 => sin_data_int <= to_signed(983,32); cos_data_int <= to_signed(-186,32);
				when 1146 => sin_data_int <= to_signed(983,32); cos_data_int <= to_signed(-188,32);
				when 1147 => sin_data_int <= to_signed(982,32); cos_data_int <= to_signed(-189,32);
				when 1148 => sin_data_int <= to_signed(982,32); cos_data_int <= to_signed(-191,32);
				when 1149 => sin_data_int <= to_signed(982,32); cos_data_int <= to_signed(-192,32);
				when 1150 => sin_data_int <= to_signed(981,32); cos_data_int <= to_signed(-194,32);
				when 1151 => sin_data_int <= to_signed(981,32); cos_data_int <= to_signed(-195,32);
				when 1152 => sin_data_int <= to_signed(981,32); cos_data_int <= to_signed(-197,32);
				when 1153 => sin_data_int <= to_signed(980,32); cos_data_int <= to_signed(-198,32);
				when 1154 => sin_data_int <= to_signed(980,32); cos_data_int <= to_signed(-200,32);
				when 1155 => sin_data_int <= to_signed(980,32); cos_data_int <= to_signed(-201,32);
				when 1156 => sin_data_int <= to_signed(980,32); cos_data_int <= to_signed(-203,32);
				when 1157 => sin_data_int <= to_signed(979,32); cos_data_int <= to_signed(-204,32);
				when 1158 => sin_data_int <= to_signed(979,32); cos_data_int <= to_signed(-206,32);
				when 1159 => sin_data_int <= to_signed(979,32); cos_data_int <= to_signed(-207,32);
				when 1160 => sin_data_int <= to_signed(978,32); cos_data_int <= to_signed(-209,32);
				when 1161 => sin_data_int <= to_signed(978,32); cos_data_int <= to_signed(-210,32);
				when 1162 => sin_data_int <= to_signed(978,32); cos_data_int <= to_signed(-212,32);
				when 1163 => sin_data_int <= to_signed(977,32); cos_data_int <= to_signed(-213,32);
				when 1164 => sin_data_int <= to_signed(977,32); cos_data_int <= to_signed(-215,32);
				when 1165 => sin_data_int <= to_signed(977,32); cos_data_int <= to_signed(-216,32);
				when 1166 => sin_data_int <= to_signed(976,32); cos_data_int <= to_signed(-218,32);
				when 1167 => sin_data_int <= to_signed(976,32); cos_data_int <= to_signed(-219,32);
				when 1168 => sin_data_int <= to_signed(976,32); cos_data_int <= to_signed(-221,32);
				when 1169 => sin_data_int <= to_signed(975,32); cos_data_int <= to_signed(-222,32);
				when 1170 => sin_data_int <= to_signed(975,32); cos_data_int <= to_signed(-224,32);
				when 1171 => sin_data_int <= to_signed(975,32); cos_data_int <= to_signed(-225,32);
				when 1172 => sin_data_int <= to_signed(974,32); cos_data_int <= to_signed(-227,32);
				when 1173 => sin_data_int <= to_signed(974,32); cos_data_int <= to_signed(-228,32);
				when 1174 => sin_data_int <= to_signed(974,32); cos_data_int <= to_signed(-230,32);
				when 1175 => sin_data_int <= to_signed(973,32); cos_data_int <= to_signed(-231,32);
				when 1176 => sin_data_int <= to_signed(973,32); cos_data_int <= to_signed(-233,32);
				when 1177 => sin_data_int <= to_signed(973,32); cos_data_int <= to_signed(-234,32);
				when 1178 => sin_data_int <= to_signed(972,32); cos_data_int <= to_signed(-236,32);
				when 1179 => sin_data_int <= to_signed(972,32); cos_data_int <= to_signed(-237,32);
				when 1180 => sin_data_int <= to_signed(972,32); cos_data_int <= to_signed(-239,32);
				when 1181 => sin_data_int <= to_signed(971,32); cos_data_int <= to_signed(-240,32);
				when 1182 => sin_data_int <= to_signed(971,32); cos_data_int <= to_signed(-241,32);
				when 1183 => sin_data_int <= to_signed(970,32); cos_data_int <= to_signed(-243,32);
				when 1184 => sin_data_int <= to_signed(970,32); cos_data_int <= to_signed(-244,32);
				when 1185 => sin_data_int <= to_signed(970,32); cos_data_int <= to_signed(-246,32);
				when 1186 => sin_data_int <= to_signed(969,32); cos_data_int <= to_signed(-247,32);
				when 1187 => sin_data_int <= to_signed(969,32); cos_data_int <= to_signed(-249,32);
				when 1188 => sin_data_int <= to_signed(969,32); cos_data_int <= to_signed(-250,32);
				when 1189 => sin_data_int <= to_signed(968,32); cos_data_int <= to_signed(-252,32);
				when 1190 => sin_data_int <= to_signed(968,32); cos_data_int <= to_signed(-253,32);
				when 1191 => sin_data_int <= to_signed(967,32); cos_data_int <= to_signed(-255,32);
				when 1192 => sin_data_int <= to_signed(967,32); cos_data_int <= to_signed(-256,32);
				when 1193 => sin_data_int <= to_signed(967,32); cos_data_int <= to_signed(-258,32);
				when 1194 => sin_data_int <= to_signed(966,32); cos_data_int <= to_signed(-259,32);
				when 1195 => sin_data_int <= to_signed(966,32); cos_data_int <= to_signed(-261,32);
				when 1196 => sin_data_int <= to_signed(965,32); cos_data_int <= to_signed(-262,32);
				when 1197 => sin_data_int <= to_signed(965,32); cos_data_int <= to_signed(-264,32);
				when 1198 => sin_data_int <= to_signed(965,32); cos_data_int <= to_signed(-265,32);
				when 1199 => sin_data_int <= to_signed(964,32); cos_data_int <= to_signed(-267,32);
				when 1200 => sin_data_int <= to_signed(964,32); cos_data_int <= to_signed(-268,32);
				when 1201 => sin_data_int <= to_signed(963,32); cos_data_int <= to_signed(-270,32);
				when 1202 => sin_data_int <= to_signed(963,32); cos_data_int <= to_signed(-271,32);
				when 1203 => sin_data_int <= to_signed(963,32); cos_data_int <= to_signed(-273,32);
				when 1204 => sin_data_int <= to_signed(962,32); cos_data_int <= to_signed(-274,32);
				when 1205 => sin_data_int <= to_signed(962,32); cos_data_int <= to_signed(-276,32);
				when 1206 => sin_data_int <= to_signed(961,32); cos_data_int <= to_signed(-277,32);
				when 1207 => sin_data_int <= to_signed(961,32); cos_data_int <= to_signed(-279,32);
				when 1208 => sin_data_int <= to_signed(960,32); cos_data_int <= to_signed(-280,32);
				when 1209 => sin_data_int <= to_signed(960,32); cos_data_int <= to_signed(-281,32);
				when 1210 => sin_data_int <= to_signed(960,32); cos_data_int <= to_signed(-283,32);
				when 1211 => sin_data_int <= to_signed(959,32); cos_data_int <= to_signed(-284,32);
				when 1212 => sin_data_int <= to_signed(959,32); cos_data_int <= to_signed(-286,32);
				when 1213 => sin_data_int <= to_signed(958,32); cos_data_int <= to_signed(-287,32);
				when 1214 => sin_data_int <= to_signed(958,32); cos_data_int <= to_signed(-289,32);
				when 1215 => sin_data_int <= to_signed(957,32); cos_data_int <= to_signed(-290,32);
				when 1216 => sin_data_int <= to_signed(957,32); cos_data_int <= to_signed(-292,32);
				when 1217 => sin_data_int <= to_signed(956,32); cos_data_int <= to_signed(-293,32);
				when 1218 => sin_data_int <= to_signed(956,32); cos_data_int <= to_signed(-295,32);
				when 1219 => sin_data_int <= to_signed(956,32); cos_data_int <= to_signed(-296,32);
				when 1220 => sin_data_int <= to_signed(955,32); cos_data_int <= to_signed(-298,32);
				when 1221 => sin_data_int <= to_signed(955,32); cos_data_int <= to_signed(-299,32);
				when 1222 => sin_data_int <= to_signed(954,32); cos_data_int <= to_signed(-301,32);
				when 1223 => sin_data_int <= to_signed(954,32); cos_data_int <= to_signed(-302,32);
				when 1224 => sin_data_int <= to_signed(953,32); cos_data_int <= to_signed(-303,32);
				when 1225 => sin_data_int <= to_signed(953,32); cos_data_int <= to_signed(-305,32);
				when 1226 => sin_data_int <= to_signed(952,32); cos_data_int <= to_signed(-306,32);
				when 1227 => sin_data_int <= to_signed(952,32); cos_data_int <= to_signed(-308,32);
				when 1228 => sin_data_int <= to_signed(951,32); cos_data_int <= to_signed(-309,32);
				when 1229 => sin_data_int <= to_signed(951,32); cos_data_int <= to_signed(-311,32);
				when 1230 => sin_data_int <= to_signed(950,32); cos_data_int <= to_signed(-312,32);
				when 1231 => sin_data_int <= to_signed(950,32); cos_data_int <= to_signed(-314,32);
				when 1232 => sin_data_int <= to_signed(950,32); cos_data_int <= to_signed(-315,32);
				when 1233 => sin_data_int <= to_signed(949,32); cos_data_int <= to_signed(-317,32);
				when 1234 => sin_data_int <= to_signed(949,32); cos_data_int <= to_signed(-318,32);
				when 1235 => sin_data_int <= to_signed(948,32); cos_data_int <= to_signed(-320,32);
				when 1236 => sin_data_int <= to_signed(948,32); cos_data_int <= to_signed(-321,32);
				when 1237 => sin_data_int <= to_signed(947,32); cos_data_int <= to_signed(-322,32);
				when 1238 => sin_data_int <= to_signed(947,32); cos_data_int <= to_signed(-324,32);
				when 1239 => sin_data_int <= to_signed(946,32); cos_data_int <= to_signed(-325,32);
				when 1240 => sin_data_int <= to_signed(946,32); cos_data_int <= to_signed(-327,32);
				when 1241 => sin_data_int <= to_signed(945,32); cos_data_int <= to_signed(-328,32);
				when 1242 => sin_data_int <= to_signed(945,32); cos_data_int <= to_signed(-330,32);
				when 1243 => sin_data_int <= to_signed(944,32); cos_data_int <= to_signed(-331,32);
				when 1244 => sin_data_int <= to_signed(944,32); cos_data_int <= to_signed(-333,32);
				when 1245 => sin_data_int <= to_signed(943,32); cos_data_int <= to_signed(-334,32);
				when 1246 => sin_data_int <= to_signed(943,32); cos_data_int <= to_signed(-335,32);
				when 1247 => sin_data_int <= to_signed(942,32); cos_data_int <= to_signed(-337,32);
				when 1248 => sin_data_int <= to_signed(942,32); cos_data_int <= to_signed(-338,32);
				when 1249 => sin_data_int <= to_signed(941,32); cos_data_int <= to_signed(-340,32);
				when 1250 => sin_data_int <= to_signed(941,32); cos_data_int <= to_signed(-341,32);
				when 1251 => sin_data_int <= to_signed(940,32); cos_data_int <= to_signed(-343,32);
				when 1252 => sin_data_int <= to_signed(939,32); cos_data_int <= to_signed(-344,32);
				when 1253 => sin_data_int <= to_signed(939,32); cos_data_int <= to_signed(-346,32);
				when 1254 => sin_data_int <= to_signed(938,32); cos_data_int <= to_signed(-347,32);
				when 1255 => sin_data_int <= to_signed(938,32); cos_data_int <= to_signed(-348,32);
				when 1256 => sin_data_int <= to_signed(937,32); cos_data_int <= to_signed(-350,32);
				when 1257 => sin_data_int <= to_signed(937,32); cos_data_int <= to_signed(-351,32);
				when 1258 => sin_data_int <= to_signed(936,32); cos_data_int <= to_signed(-353,32);
				when 1259 => sin_data_int <= to_signed(936,32); cos_data_int <= to_signed(-354,32);
				when 1260 => sin_data_int <= to_signed(935,32); cos_data_int <= to_signed(-356,32);
				when 1261 => sin_data_int <= to_signed(935,32); cos_data_int <= to_signed(-357,32);
				when 1262 => sin_data_int <= to_signed(934,32); cos_data_int <= to_signed(-358,32);
				when 1263 => sin_data_int <= to_signed(934,32); cos_data_int <= to_signed(-360,32);
				when 1264 => sin_data_int <= to_signed(933,32); cos_data_int <= to_signed(-361,32);
				when 1265 => sin_data_int <= to_signed(932,32); cos_data_int <= to_signed(-363,32);
				when 1266 => sin_data_int <= to_signed(932,32); cos_data_int <= to_signed(-364,32);
				when 1267 => sin_data_int <= to_signed(931,32); cos_data_int <= to_signed(-366,32);
				when 1268 => sin_data_int <= to_signed(931,32); cos_data_int <= to_signed(-367,32);
				when 1269 => sin_data_int <= to_signed(930,32); cos_data_int <= to_signed(-368,32);
				when 1270 => sin_data_int <= to_signed(930,32); cos_data_int <= to_signed(-370,32);
				when 1271 => sin_data_int <= to_signed(929,32); cos_data_int <= to_signed(-371,32);
				when 1272 => sin_data_int <= to_signed(929,32); cos_data_int <= to_signed(-373,32);
				when 1273 => sin_data_int <= to_signed(928,32); cos_data_int <= to_signed(-374,32);
				when 1274 => sin_data_int <= to_signed(927,32); cos_data_int <= to_signed(-376,32);
				when 1275 => sin_data_int <= to_signed(927,32); cos_data_int <= to_signed(-377,32);
				when 1276 => sin_data_int <= to_signed(926,32); cos_data_int <= to_signed(-378,32);
				when 1277 => sin_data_int <= to_signed(926,32); cos_data_int <= to_signed(-380,32);
				when 1278 => sin_data_int <= to_signed(925,32); cos_data_int <= to_signed(-381,32);
				when 1279 => sin_data_int <= to_signed(924,32); cos_data_int <= to_signed(-383,32);
				when 1280 => sin_data_int <= to_signed(924,32); cos_data_int <= to_signed(-384,32);
				when 1281 => sin_data_int <= to_signed(923,32); cos_data_int <= to_signed(-386,32);
				when 1282 => sin_data_int <= to_signed(923,32); cos_data_int <= to_signed(-387,32);
				when 1283 => sin_data_int <= to_signed(922,32); cos_data_int <= to_signed(-388,32);
				when 1284 => sin_data_int <= to_signed(922,32); cos_data_int <= to_signed(-390,32);
				when 1285 => sin_data_int <= to_signed(921,32); cos_data_int <= to_signed(-391,32);
				when 1286 => sin_data_int <= to_signed(920,32); cos_data_int <= to_signed(-393,32);
				when 1287 => sin_data_int <= to_signed(920,32); cos_data_int <= to_signed(-394,32);
				when 1288 => sin_data_int <= to_signed(919,32); cos_data_int <= to_signed(-395,32);
				when 1289 => sin_data_int <= to_signed(919,32); cos_data_int <= to_signed(-397,32);
				when 1290 => sin_data_int <= to_signed(918,32); cos_data_int <= to_signed(-398,32);
				when 1291 => sin_data_int <= to_signed(917,32); cos_data_int <= to_signed(-400,32);
				when 1292 => sin_data_int <= to_signed(917,32); cos_data_int <= to_signed(-401,32);
				when 1293 => sin_data_int <= to_signed(916,32); cos_data_int <= to_signed(-402,32);
				when 1294 => sin_data_int <= to_signed(915,32); cos_data_int <= to_signed(-404,32);
				when 1295 => sin_data_int <= to_signed(915,32); cos_data_int <= to_signed(-405,32);
				when 1296 => sin_data_int <= to_signed(914,32); cos_data_int <= to_signed(-407,32);
				when 1297 => sin_data_int <= to_signed(914,32); cos_data_int <= to_signed(-408,32);
				when 1298 => sin_data_int <= to_signed(913,32); cos_data_int <= to_signed(-409,32);
				when 1299 => sin_data_int <= to_signed(912,32); cos_data_int <= to_signed(-411,32);
				when 1300 => sin_data_int <= to_signed(912,32); cos_data_int <= to_signed(-412,32);
				when 1301 => sin_data_int <= to_signed(911,32); cos_data_int <= to_signed(-414,32);
				when 1302 => sin_data_int <= to_signed(910,32); cos_data_int <= to_signed(-415,32);
				when 1303 => sin_data_int <= to_signed(910,32); cos_data_int <= to_signed(-416,32);
				when 1304 => sin_data_int <= to_signed(909,32); cos_data_int <= to_signed(-418,32);
				when 1305 => sin_data_int <= to_signed(909,32); cos_data_int <= to_signed(-419,32);
				when 1306 => sin_data_int <= to_signed(908,32); cos_data_int <= to_signed(-421,32);
				when 1307 => sin_data_int <= to_signed(907,32); cos_data_int <= to_signed(-422,32);
				when 1308 => sin_data_int <= to_signed(907,32); cos_data_int <= to_signed(-423,32);
				when 1309 => sin_data_int <= to_signed(906,32); cos_data_int <= to_signed(-425,32);
				when 1310 => sin_data_int <= to_signed(905,32); cos_data_int <= to_signed(-426,32);
				when 1311 => sin_data_int <= to_signed(905,32); cos_data_int <= to_signed(-428,32);
				when 1312 => sin_data_int <= to_signed(904,32); cos_data_int <= to_signed(-429,32);
				when 1313 => sin_data_int <= to_signed(903,32); cos_data_int <= to_signed(-430,32);
				when 1314 => sin_data_int <= to_signed(903,32); cos_data_int <= to_signed(-432,32);
				when 1315 => sin_data_int <= to_signed(902,32); cos_data_int <= to_signed(-433,32);
				when 1316 => sin_data_int <= to_signed(901,32); cos_data_int <= to_signed(-434,32);
				when 1317 => sin_data_int <= to_signed(901,32); cos_data_int <= to_signed(-436,32);
				when 1318 => sin_data_int <= to_signed(900,32); cos_data_int <= to_signed(-437,32);
				when 1319 => sin_data_int <= to_signed(899,32); cos_data_int <= to_signed(-439,32);
				when 1320 => sin_data_int <= to_signed(899,32); cos_data_int <= to_signed(-440,32);
				when 1321 => sin_data_int <= to_signed(898,32); cos_data_int <= to_signed(-441,32);
				when 1322 => sin_data_int <= to_signed(897,32); cos_data_int <= to_signed(-443,32);
				when 1323 => sin_data_int <= to_signed(897,32); cos_data_int <= to_signed(-444,32);
				when 1324 => sin_data_int <= to_signed(896,32); cos_data_int <= to_signed(-445,32);
				when 1325 => sin_data_int <= to_signed(895,32); cos_data_int <= to_signed(-447,32);
				when 1326 => sin_data_int <= to_signed(895,32); cos_data_int <= to_signed(-448,32);
				when 1327 => sin_data_int <= to_signed(894,32); cos_data_int <= to_signed(-450,32);
				when 1328 => sin_data_int <= to_signed(893,32); cos_data_int <= to_signed(-451,32);
				when 1329 => sin_data_int <= to_signed(893,32); cos_data_int <= to_signed(-452,32);
				when 1330 => sin_data_int <= to_signed(892,32); cos_data_int <= to_signed(-454,32);
				when 1331 => sin_data_int <= to_signed(891,32); cos_data_int <= to_signed(-455,32);
				when 1332 => sin_data_int <= to_signed(890,32); cos_data_int <= to_signed(-456,32);
				when 1333 => sin_data_int <= to_signed(890,32); cos_data_int <= to_signed(-458,32);
				when 1334 => sin_data_int <= to_signed(889,32); cos_data_int <= to_signed(-459,32);
				when 1335 => sin_data_int <= to_signed(888,32); cos_data_int <= to_signed(-461,32);
				when 1336 => sin_data_int <= to_signed(888,32); cos_data_int <= to_signed(-462,32);
				when 1337 => sin_data_int <= to_signed(887,32); cos_data_int <= to_signed(-463,32);
				when 1338 => sin_data_int <= to_signed(886,32); cos_data_int <= to_signed(-465,32);
				when 1339 => sin_data_int <= to_signed(886,32); cos_data_int <= to_signed(-466,32);
				when 1340 => sin_data_int <= to_signed(885,32); cos_data_int <= to_signed(-467,32);
				when 1341 => sin_data_int <= to_signed(884,32); cos_data_int <= to_signed(-469,32);
				when 1342 => sin_data_int <= to_signed(883,32); cos_data_int <= to_signed(-470,32);
				when 1343 => sin_data_int <= to_signed(883,32); cos_data_int <= to_signed(-471,32);
				when 1344 => sin_data_int <= to_signed(882,32); cos_data_int <= to_signed(-473,32);
				when 1345 => sin_data_int <= to_signed(881,32); cos_data_int <= to_signed(-474,32);
				when 1346 => sin_data_int <= to_signed(880,32); cos_data_int <= to_signed(-475,32);
				when 1347 => sin_data_int <= to_signed(880,32); cos_data_int <= to_signed(-477,32);
				when 1348 => sin_data_int <= to_signed(879,32); cos_data_int <= to_signed(-478,32);
				when 1349 => sin_data_int <= to_signed(878,32); cos_data_int <= to_signed(-479,32);
				when 1350 => sin_data_int <= to_signed(878,32); cos_data_int <= to_signed(-481,32);
				when 1351 => sin_data_int <= to_signed(877,32); cos_data_int <= to_signed(-482,32);
				when 1352 => sin_data_int <= to_signed(876,32); cos_data_int <= to_signed(-484,32);
				when 1353 => sin_data_int <= to_signed(875,32); cos_data_int <= to_signed(-485,32);
				when 1354 => sin_data_int <= to_signed(875,32); cos_data_int <= to_signed(-486,32);
				when 1355 => sin_data_int <= to_signed(874,32); cos_data_int <= to_signed(-488,32);
				when 1356 => sin_data_int <= to_signed(873,32); cos_data_int <= to_signed(-489,32);
				when 1357 => sin_data_int <= to_signed(872,32); cos_data_int <= to_signed(-490,32);
				when 1358 => sin_data_int <= to_signed(872,32); cos_data_int <= to_signed(-492,32);
				when 1359 => sin_data_int <= to_signed(871,32); cos_data_int <= to_signed(-493,32);
				when 1360 => sin_data_int <= to_signed(870,32); cos_data_int <= to_signed(-494,32);
				when 1361 => sin_data_int <= to_signed(869,32); cos_data_int <= to_signed(-496,32);
				when 1362 => sin_data_int <= to_signed(869,32); cos_data_int <= to_signed(-497,32);
				when 1363 => sin_data_int <= to_signed(868,32); cos_data_int <= to_signed(-498,32);
				when 1364 => sin_data_int <= to_signed(867,32); cos_data_int <= to_signed(-500,32);
				when 1365 => sin_data_int <= to_signed(866,32); cos_data_int <= to_signed(-501,32);
				when 1366 => sin_data_int <= to_signed(866,32); cos_data_int <= to_signed(-502,32);
				when 1367 => sin_data_int <= to_signed(865,32); cos_data_int <= to_signed(-504,32);
				when 1368 => sin_data_int <= to_signed(864,32); cos_data_int <= to_signed(-505,32);
				when 1369 => sin_data_int <= to_signed(863,32); cos_data_int <= to_signed(-506,32);
				when 1370 => sin_data_int <= to_signed(862,32); cos_data_int <= to_signed(-508,32);
				when 1371 => sin_data_int <= to_signed(862,32); cos_data_int <= to_signed(-509,32);
				when 1372 => sin_data_int <= to_signed(861,32); cos_data_int <= to_signed(-510,32);
				when 1373 => sin_data_int <= to_signed(860,32); cos_data_int <= to_signed(-511,32);
				when 1374 => sin_data_int <= to_signed(859,32); cos_data_int <= to_signed(-513,32);
				when 1375 => sin_data_int <= to_signed(859,32); cos_data_int <= to_signed(-514,32);
				when 1376 => sin_data_int <= to_signed(858,32); cos_data_int <= to_signed(-515,32);
				when 1377 => sin_data_int <= to_signed(857,32); cos_data_int <= to_signed(-517,32);
				when 1378 => sin_data_int <= to_signed(856,32); cos_data_int <= to_signed(-518,32);
				when 1379 => sin_data_int <= to_signed(855,32); cos_data_int <= to_signed(-519,32);
				when 1380 => sin_data_int <= to_signed(855,32); cos_data_int <= to_signed(-521,32);
				when 1381 => sin_data_int <= to_signed(854,32); cos_data_int <= to_signed(-522,32);
				when 1382 => sin_data_int <= to_signed(853,32); cos_data_int <= to_signed(-523,32);
				when 1383 => sin_data_int <= to_signed(852,32); cos_data_int <= to_signed(-525,32);
				when 1384 => sin_data_int <= to_signed(851,32); cos_data_int <= to_signed(-526,32);
				when 1385 => sin_data_int <= to_signed(851,32); cos_data_int <= to_signed(-527,32);
				when 1386 => sin_data_int <= to_signed(850,32); cos_data_int <= to_signed(-529,32);
				when 1387 => sin_data_int <= to_signed(849,32); cos_data_int <= to_signed(-530,32);
				when 1388 => sin_data_int <= to_signed(848,32); cos_data_int <= to_signed(-531,32);
				when 1389 => sin_data_int <= to_signed(847,32); cos_data_int <= to_signed(-532,32);
				when 1390 => sin_data_int <= to_signed(846,32); cos_data_int <= to_signed(-534,32);
				when 1391 => sin_data_int <= to_signed(846,32); cos_data_int <= to_signed(-535,32);
				when 1392 => sin_data_int <= to_signed(845,32); cos_data_int <= to_signed(-536,32);
				when 1393 => sin_data_int <= to_signed(844,32); cos_data_int <= to_signed(-538,32);
				when 1394 => sin_data_int <= to_signed(843,32); cos_data_int <= to_signed(-539,32);
				when 1395 => sin_data_int <= to_signed(842,32); cos_data_int <= to_signed(-540,32);
				when 1396 => sin_data_int <= to_signed(842,32); cos_data_int <= to_signed(-541,32);
				when 1397 => sin_data_int <= to_signed(841,32); cos_data_int <= to_signed(-543,32);
				when 1398 => sin_data_int <= to_signed(840,32); cos_data_int <= to_signed(-544,32);
				when 1399 => sin_data_int <= to_signed(839,32); cos_data_int <= to_signed(-545,32);
				when 1400 => sin_data_int <= to_signed(838,32); cos_data_int <= to_signed(-547,32);
				when 1401 => sin_data_int <= to_signed(837,32); cos_data_int <= to_signed(-548,32);
				when 1402 => sin_data_int <= to_signed(837,32); cos_data_int <= to_signed(-549,32);
				when 1403 => sin_data_int <= to_signed(836,32); cos_data_int <= to_signed(-550,32);
				when 1404 => sin_data_int <= to_signed(835,32); cos_data_int <= to_signed(-552,32);
				when 1405 => sin_data_int <= to_signed(834,32); cos_data_int <= to_signed(-553,32);
				when 1406 => sin_data_int <= to_signed(833,32); cos_data_int <= to_signed(-554,32);
				when 1407 => sin_data_int <= to_signed(832,32); cos_data_int <= to_signed(-556,32);
				when 1408 => sin_data_int <= to_signed(831,32); cos_data_int <= to_signed(-557,32);
				when 1409 => sin_data_int <= to_signed(831,32); cos_data_int <= to_signed(-558,32);
				when 1410 => sin_data_int <= to_signed(830,32); cos_data_int <= to_signed(-559,32);
				when 1411 => sin_data_int <= to_signed(829,32); cos_data_int <= to_signed(-561,32);
				when 1412 => sin_data_int <= to_signed(828,32); cos_data_int <= to_signed(-562,32);
				when 1413 => sin_data_int <= to_signed(827,32); cos_data_int <= to_signed(-563,32);
				when 1414 => sin_data_int <= to_signed(826,32); cos_data_int <= to_signed(-564,32);
				when 1415 => sin_data_int <= to_signed(825,32); cos_data_int <= to_signed(-566,32);
				when 1416 => sin_data_int <= to_signed(825,32); cos_data_int <= to_signed(-567,32);
				when 1417 => sin_data_int <= to_signed(824,32); cos_data_int <= to_signed(-568,32);
				when 1418 => sin_data_int <= to_signed(823,32); cos_data_int <= to_signed(-570,32);
				when 1419 => sin_data_int <= to_signed(822,32); cos_data_int <= to_signed(-571,32);
				when 1420 => sin_data_int <= to_signed(821,32); cos_data_int <= to_signed(-572,32);
				when 1421 => sin_data_int <= to_signed(820,32); cos_data_int <= to_signed(-573,32);
				when 1422 => sin_data_int <= to_signed(819,32); cos_data_int <= to_signed(-575,32);
				when 1423 => sin_data_int <= to_signed(818,32); cos_data_int <= to_signed(-576,32);
				when 1424 => sin_data_int <= to_signed(818,32); cos_data_int <= to_signed(-577,32);
				when 1425 => sin_data_int <= to_signed(817,32); cos_data_int <= to_signed(-578,32);
				when 1426 => sin_data_int <= to_signed(816,32); cos_data_int <= to_signed(-580,32);
				when 1427 => sin_data_int <= to_signed(815,32); cos_data_int <= to_signed(-581,32);
				when 1428 => sin_data_int <= to_signed(814,32); cos_data_int <= to_signed(-582,32);
				when 1429 => sin_data_int <= to_signed(813,32); cos_data_int <= to_signed(-583,32);
				when 1430 => sin_data_int <= to_signed(812,32); cos_data_int <= to_signed(-585,32);
				when 1431 => sin_data_int <= to_signed(811,32); cos_data_int <= to_signed(-586,32);
				when 1432 => sin_data_int <= to_signed(810,32); cos_data_int <= to_signed(-587,32);
				when 1433 => sin_data_int <= to_signed(810,32); cos_data_int <= to_signed(-588,32);
				when 1434 => sin_data_int <= to_signed(809,32); cos_data_int <= to_signed(-590,32);
				when 1435 => sin_data_int <= to_signed(808,32); cos_data_int <= to_signed(-591,32);
				when 1436 => sin_data_int <= to_signed(807,32); cos_data_int <= to_signed(-592,32);
				when 1437 => sin_data_int <= to_signed(806,32); cos_data_int <= to_signed(-593,32);
				when 1438 => sin_data_int <= to_signed(805,32); cos_data_int <= to_signed(-594,32);
				when 1439 => sin_data_int <= to_signed(804,32); cos_data_int <= to_signed(-596,32);
				when 1440 => sin_data_int <= to_signed(803,32); cos_data_int <= to_signed(-597,32);
				when 1441 => sin_data_int <= to_signed(802,32); cos_data_int <= to_signed(-598,32);
				when 1442 => sin_data_int <= to_signed(801,32); cos_data_int <= to_signed(-599,32);
				when 1443 => sin_data_int <= to_signed(800,32); cos_data_int <= to_signed(-601,32);
				when 1444 => sin_data_int <= to_signed(800,32); cos_data_int <= to_signed(-602,32);
				when 1445 => sin_data_int <= to_signed(799,32); cos_data_int <= to_signed(-603,32);
				when 1446 => sin_data_int <= to_signed(798,32); cos_data_int <= to_signed(-604,32);
				when 1447 => sin_data_int <= to_signed(797,32); cos_data_int <= to_signed(-606,32);
				when 1448 => sin_data_int <= to_signed(796,32); cos_data_int <= to_signed(-607,32);
				when 1449 => sin_data_int <= to_signed(795,32); cos_data_int <= to_signed(-608,32);
				when 1450 => sin_data_int <= to_signed(794,32); cos_data_int <= to_signed(-609,32);
				when 1451 => sin_data_int <= to_signed(793,32); cos_data_int <= to_signed(-610,32);
				when 1452 => sin_data_int <= to_signed(792,32); cos_data_int <= to_signed(-612,32);
				when 1453 => sin_data_int <= to_signed(791,32); cos_data_int <= to_signed(-613,32);
				when 1454 => sin_data_int <= to_signed(790,32); cos_data_int <= to_signed(-614,32);
				when 1455 => sin_data_int <= to_signed(789,32); cos_data_int <= to_signed(-615,32);
				when 1456 => sin_data_int <= to_signed(788,32); cos_data_int <= to_signed(-616,32);
				when 1457 => sin_data_int <= to_signed(787,32); cos_data_int <= to_signed(-618,32);
				when 1458 => sin_data_int <= to_signed(786,32); cos_data_int <= to_signed(-619,32);
				when 1459 => sin_data_int <= to_signed(786,32); cos_data_int <= to_signed(-620,32);
				when 1460 => sin_data_int <= to_signed(785,32); cos_data_int <= to_signed(-621,32);
				when 1461 => sin_data_int <= to_signed(784,32); cos_data_int <= to_signed(-622,32);
				when 1462 => sin_data_int <= to_signed(783,32); cos_data_int <= to_signed(-624,32);
				when 1463 => sin_data_int <= to_signed(782,32); cos_data_int <= to_signed(-625,32);
				when 1464 => sin_data_int <= to_signed(781,32); cos_data_int <= to_signed(-626,32);
				when 1465 => sin_data_int <= to_signed(780,32); cos_data_int <= to_signed(-627,32);
				when 1466 => sin_data_int <= to_signed(779,32); cos_data_int <= to_signed(-628,32);
				when 1467 => sin_data_int <= to_signed(778,32); cos_data_int <= to_signed(-630,32);
				when 1468 => sin_data_int <= to_signed(777,32); cos_data_int <= to_signed(-631,32);
				when 1469 => sin_data_int <= to_signed(776,32); cos_data_int <= to_signed(-632,32);
				when 1470 => sin_data_int <= to_signed(775,32); cos_data_int <= to_signed(-633,32);
				when 1471 => sin_data_int <= to_signed(774,32); cos_data_int <= to_signed(-634,32);
				when 1472 => sin_data_int <= to_signed(773,32); cos_data_int <= to_signed(-636,32);
				when 1473 => sin_data_int <= to_signed(772,32); cos_data_int <= to_signed(-637,32);
				when 1474 => sin_data_int <= to_signed(771,32); cos_data_int <= to_signed(-638,32);
				when 1475 => sin_data_int <= to_signed(770,32); cos_data_int <= to_signed(-639,32);
				when 1476 => sin_data_int <= to_signed(769,32); cos_data_int <= to_signed(-640,32);
				when 1477 => sin_data_int <= to_signed(768,32); cos_data_int <= to_signed(-641,32);
				when 1478 => sin_data_int <= to_signed(767,32); cos_data_int <= to_signed(-643,32);
				when 1479 => sin_data_int <= to_signed(766,32); cos_data_int <= to_signed(-644,32);
				when 1480 => sin_data_int <= to_signed(765,32); cos_data_int <= to_signed(-645,32);
				when 1481 => sin_data_int <= to_signed(764,32); cos_data_int <= to_signed(-646,32);
				when 1482 => sin_data_int <= to_signed(763,32); cos_data_int <= to_signed(-647,32);
				when 1483 => sin_data_int <= to_signed(762,32); cos_data_int <= to_signed(-649,32);
				when 1484 => sin_data_int <= to_signed(761,32); cos_data_int <= to_signed(-650,32);
				when 1485 => sin_data_int <= to_signed(760,32); cos_data_int <= to_signed(-651,32);
				when 1486 => sin_data_int <= to_signed(759,32); cos_data_int <= to_signed(-652,32);
				when 1487 => sin_data_int <= to_signed(758,32); cos_data_int <= to_signed(-653,32);
				when 1488 => sin_data_int <= to_signed(757,32); cos_data_int <= to_signed(-654,32);
				when 1489 => sin_data_int <= to_signed(756,32); cos_data_int <= to_signed(-655,32);
				when 1490 => sin_data_int <= to_signed(755,32); cos_data_int <= to_signed(-657,32);
				when 1491 => sin_data_int <= to_signed(754,32); cos_data_int <= to_signed(-658,32);
				when 1492 => sin_data_int <= to_signed(753,32); cos_data_int <= to_signed(-659,32);
				when 1493 => sin_data_int <= to_signed(752,32); cos_data_int <= to_signed(-660,32);
				when 1494 => sin_data_int <= to_signed(751,32); cos_data_int <= to_signed(-661,32);
				when 1495 => sin_data_int <= to_signed(750,32); cos_data_int <= to_signed(-662,32);
				when 1496 => sin_data_int <= to_signed(749,32); cos_data_int <= to_signed(-664,32);
				when 1497 => sin_data_int <= to_signed(748,32); cos_data_int <= to_signed(-665,32);
				when 1498 => sin_data_int <= to_signed(747,32); cos_data_int <= to_signed(-666,32);
				when 1499 => sin_data_int <= to_signed(746,32); cos_data_int <= to_signed(-667,32);
				when 1500 => sin_data_int <= to_signed(745,32); cos_data_int <= to_signed(-668,32);
				when 1501 => sin_data_int <= to_signed(744,32); cos_data_int <= to_signed(-669,32);
				when 1502 => sin_data_int <= to_signed(743,32); cos_data_int <= to_signed(-670,32);
				when 1503 => sin_data_int <= to_signed(742,32); cos_data_int <= to_signed(-672,32);
				when 1504 => sin_data_int <= to_signed(741,32); cos_data_int <= to_signed(-673,32);
				when 1505 => sin_data_int <= to_signed(740,32); cos_data_int <= to_signed(-674,32);
				when 1506 => sin_data_int <= to_signed(739,32); cos_data_int <= to_signed(-675,32);
				when 1507 => sin_data_int <= to_signed(738,32); cos_data_int <= to_signed(-676,32);
				when 1508 => sin_data_int <= to_signed(737,32); cos_data_int <= to_signed(-677,32);
				when 1509 => sin_data_int <= to_signed(736,32); cos_data_int <= to_signed(-678,32);
				when 1510 => sin_data_int <= to_signed(735,32); cos_data_int <= to_signed(-679,32);
				when 1511 => sin_data_int <= to_signed(734,32); cos_data_int <= to_signed(-681,32);
				when 1512 => sin_data_int <= to_signed(733,32); cos_data_int <= to_signed(-682,32);
				when 1513 => sin_data_int <= to_signed(732,32); cos_data_int <= to_signed(-683,32);
				when 1514 => sin_data_int <= to_signed(731,32); cos_data_int <= to_signed(-684,32);
				when 1515 => sin_data_int <= to_signed(730,32); cos_data_int <= to_signed(-685,32);
				when 1516 => sin_data_int <= to_signed(728,32); cos_data_int <= to_signed(-686,32);
				when 1517 => sin_data_int <= to_signed(727,32); cos_data_int <= to_signed(-687,32);
				when 1518 => sin_data_int <= to_signed(726,32); cos_data_int <= to_signed(-688,32);
				when 1519 => sin_data_int <= to_signed(725,32); cos_data_int <= to_signed(-690,32);
				when 1520 => sin_data_int <= to_signed(724,32); cos_data_int <= to_signed(-691,32);
				when 1521 => sin_data_int <= to_signed(723,32); cos_data_int <= to_signed(-692,32);
				when 1522 => sin_data_int <= to_signed(722,32); cos_data_int <= to_signed(-693,32);
				when 1523 => sin_data_int <= to_signed(721,32); cos_data_int <= to_signed(-694,32);
				when 1524 => sin_data_int <= to_signed(720,32); cos_data_int <= to_signed(-695,32);
				when 1525 => sin_data_int <= to_signed(719,32); cos_data_int <= to_signed(-696,32);
				when 1526 => sin_data_int <= to_signed(718,32); cos_data_int <= to_signed(-697,32);
				when 1527 => sin_data_int <= to_signed(717,32); cos_data_int <= to_signed(-698,32);
				when 1528 => sin_data_int <= to_signed(716,32); cos_data_int <= to_signed(-699,32);
				when 1529 => sin_data_int <= to_signed(715,32); cos_data_int <= to_signed(-701,32);
				when 1530 => sin_data_int <= to_signed(714,32); cos_data_int <= to_signed(-702,32);
				when 1531 => sin_data_int <= to_signed(713,32); cos_data_int <= to_signed(-703,32);
				when 1532 => sin_data_int <= to_signed(711,32); cos_data_int <= to_signed(-704,32);
				when 1533 => sin_data_int <= to_signed(710,32); cos_data_int <= to_signed(-705,32);
				when 1534 => sin_data_int <= to_signed(709,32); cos_data_int <= to_signed(-706,32);
				when 1535 => sin_data_int <= to_signed(708,32); cos_data_int <= to_signed(-707,32);
				when 1536 => sin_data_int <= to_signed(707,32); cos_data_int <= to_signed(-708,32);
				when 1537 => sin_data_int <= to_signed(706,32); cos_data_int <= to_signed(-709,32);
				when 1538 => sin_data_int <= to_signed(705,32); cos_data_int <= to_signed(-710,32);
				when 1539 => sin_data_int <= to_signed(704,32); cos_data_int <= to_signed(-711,32);
				when 1540 => sin_data_int <= to_signed(703,32); cos_data_int <= to_signed(-713,32);
				when 1541 => sin_data_int <= to_signed(702,32); cos_data_int <= to_signed(-714,32);
				when 1542 => sin_data_int <= to_signed(701,32); cos_data_int <= to_signed(-715,32);
				when 1543 => sin_data_int <= to_signed(699,32); cos_data_int <= to_signed(-716,32);
				when 1544 => sin_data_int <= to_signed(698,32); cos_data_int <= to_signed(-717,32);
				when 1545 => sin_data_int <= to_signed(697,32); cos_data_int <= to_signed(-718,32);
				when 1546 => sin_data_int <= to_signed(696,32); cos_data_int <= to_signed(-719,32);
				when 1547 => sin_data_int <= to_signed(695,32); cos_data_int <= to_signed(-720,32);
				when 1548 => sin_data_int <= to_signed(694,32); cos_data_int <= to_signed(-721,32);
				when 1549 => sin_data_int <= to_signed(693,32); cos_data_int <= to_signed(-722,32);
				when 1550 => sin_data_int <= to_signed(692,32); cos_data_int <= to_signed(-723,32);
				when 1551 => sin_data_int <= to_signed(691,32); cos_data_int <= to_signed(-724,32);
				when 1552 => sin_data_int <= to_signed(690,32); cos_data_int <= to_signed(-725,32);
				when 1553 => sin_data_int <= to_signed(688,32); cos_data_int <= to_signed(-726,32);
				when 1554 => sin_data_int <= to_signed(687,32); cos_data_int <= to_signed(-727,32);
				when 1555 => sin_data_int <= to_signed(686,32); cos_data_int <= to_signed(-728,32);
				when 1556 => sin_data_int <= to_signed(685,32); cos_data_int <= to_signed(-730,32);
				when 1557 => sin_data_int <= to_signed(684,32); cos_data_int <= to_signed(-731,32);
				when 1558 => sin_data_int <= to_signed(683,32); cos_data_int <= to_signed(-732,32);
				when 1559 => sin_data_int <= to_signed(682,32); cos_data_int <= to_signed(-733,32);
				when 1560 => sin_data_int <= to_signed(681,32); cos_data_int <= to_signed(-734,32);
				when 1561 => sin_data_int <= to_signed(679,32); cos_data_int <= to_signed(-735,32);
				when 1562 => sin_data_int <= to_signed(678,32); cos_data_int <= to_signed(-736,32);
				when 1563 => sin_data_int <= to_signed(677,32); cos_data_int <= to_signed(-737,32);
				when 1564 => sin_data_int <= to_signed(676,32); cos_data_int <= to_signed(-738,32);
				when 1565 => sin_data_int <= to_signed(675,32); cos_data_int <= to_signed(-739,32);
				when 1566 => sin_data_int <= to_signed(674,32); cos_data_int <= to_signed(-740,32);
				when 1567 => sin_data_int <= to_signed(673,32); cos_data_int <= to_signed(-741,32);
				when 1568 => sin_data_int <= to_signed(672,32); cos_data_int <= to_signed(-742,32);
				when 1569 => sin_data_int <= to_signed(670,32); cos_data_int <= to_signed(-743,32);
				when 1570 => sin_data_int <= to_signed(669,32); cos_data_int <= to_signed(-744,32);
				when 1571 => sin_data_int <= to_signed(668,32); cos_data_int <= to_signed(-745,32);
				when 1572 => sin_data_int <= to_signed(667,32); cos_data_int <= to_signed(-746,32);
				when 1573 => sin_data_int <= to_signed(666,32); cos_data_int <= to_signed(-747,32);
				when 1574 => sin_data_int <= to_signed(665,32); cos_data_int <= to_signed(-748,32);
				when 1575 => sin_data_int <= to_signed(664,32); cos_data_int <= to_signed(-749,32);
				when 1576 => sin_data_int <= to_signed(662,32); cos_data_int <= to_signed(-750,32);
				when 1577 => sin_data_int <= to_signed(661,32); cos_data_int <= to_signed(-751,32);
				when 1578 => sin_data_int <= to_signed(660,32); cos_data_int <= to_signed(-752,32);
				when 1579 => sin_data_int <= to_signed(659,32); cos_data_int <= to_signed(-753,32);
				when 1580 => sin_data_int <= to_signed(658,32); cos_data_int <= to_signed(-754,32);
				when 1581 => sin_data_int <= to_signed(657,32); cos_data_int <= to_signed(-755,32);
				when 1582 => sin_data_int <= to_signed(655,32); cos_data_int <= to_signed(-756,32);
				when 1583 => sin_data_int <= to_signed(654,32); cos_data_int <= to_signed(-757,32);
				when 1584 => sin_data_int <= to_signed(653,32); cos_data_int <= to_signed(-758,32);
				when 1585 => sin_data_int <= to_signed(652,32); cos_data_int <= to_signed(-759,32);
				when 1586 => sin_data_int <= to_signed(651,32); cos_data_int <= to_signed(-760,32);
				when 1587 => sin_data_int <= to_signed(650,32); cos_data_int <= to_signed(-761,32);
				when 1588 => sin_data_int <= to_signed(649,32); cos_data_int <= to_signed(-762,32);
				when 1589 => sin_data_int <= to_signed(647,32); cos_data_int <= to_signed(-763,32);
				when 1590 => sin_data_int <= to_signed(646,32); cos_data_int <= to_signed(-764,32);
				when 1591 => sin_data_int <= to_signed(645,32); cos_data_int <= to_signed(-765,32);
				when 1592 => sin_data_int <= to_signed(644,32); cos_data_int <= to_signed(-766,32);
				when 1593 => sin_data_int <= to_signed(643,32); cos_data_int <= to_signed(-767,32);
				when 1594 => sin_data_int <= to_signed(641,32); cos_data_int <= to_signed(-768,32);
				when 1595 => sin_data_int <= to_signed(640,32); cos_data_int <= to_signed(-769,32);
				when 1596 => sin_data_int <= to_signed(639,32); cos_data_int <= to_signed(-770,32);
				when 1597 => sin_data_int <= to_signed(638,32); cos_data_int <= to_signed(-771,32);
				when 1598 => sin_data_int <= to_signed(637,32); cos_data_int <= to_signed(-772,32);
				when 1599 => sin_data_int <= to_signed(636,32); cos_data_int <= to_signed(-773,32);
				when 1600 => sin_data_int <= to_signed(634,32); cos_data_int <= to_signed(-774,32);
				when 1601 => sin_data_int <= to_signed(633,32); cos_data_int <= to_signed(-775,32);
				when 1602 => sin_data_int <= to_signed(632,32); cos_data_int <= to_signed(-776,32);
				when 1603 => sin_data_int <= to_signed(631,32); cos_data_int <= to_signed(-777,32);
				when 1604 => sin_data_int <= to_signed(630,32); cos_data_int <= to_signed(-778,32);
				when 1605 => sin_data_int <= to_signed(628,32); cos_data_int <= to_signed(-779,32);
				when 1606 => sin_data_int <= to_signed(627,32); cos_data_int <= to_signed(-780,32);
				when 1607 => sin_data_int <= to_signed(626,32); cos_data_int <= to_signed(-781,32);
				when 1608 => sin_data_int <= to_signed(625,32); cos_data_int <= to_signed(-782,32);
				when 1609 => sin_data_int <= to_signed(624,32); cos_data_int <= to_signed(-783,32);
				when 1610 => sin_data_int <= to_signed(622,32); cos_data_int <= to_signed(-784,32);
				when 1611 => sin_data_int <= to_signed(621,32); cos_data_int <= to_signed(-785,32);
				when 1612 => sin_data_int <= to_signed(620,32); cos_data_int <= to_signed(-786,32);
				when 1613 => sin_data_int <= to_signed(619,32); cos_data_int <= to_signed(-786,32);
				when 1614 => sin_data_int <= to_signed(618,32); cos_data_int <= to_signed(-787,32);
				when 1615 => sin_data_int <= to_signed(616,32); cos_data_int <= to_signed(-788,32);
				when 1616 => sin_data_int <= to_signed(615,32); cos_data_int <= to_signed(-789,32);
				when 1617 => sin_data_int <= to_signed(614,32); cos_data_int <= to_signed(-790,32);
				when 1618 => sin_data_int <= to_signed(613,32); cos_data_int <= to_signed(-791,32);
				when 1619 => sin_data_int <= to_signed(612,32); cos_data_int <= to_signed(-792,32);
				when 1620 => sin_data_int <= to_signed(610,32); cos_data_int <= to_signed(-793,32);
				when 1621 => sin_data_int <= to_signed(609,32); cos_data_int <= to_signed(-794,32);
				when 1622 => sin_data_int <= to_signed(608,32); cos_data_int <= to_signed(-795,32);
				when 1623 => sin_data_int <= to_signed(607,32); cos_data_int <= to_signed(-796,32);
				when 1624 => sin_data_int <= to_signed(606,32); cos_data_int <= to_signed(-797,32);
				when 1625 => sin_data_int <= to_signed(604,32); cos_data_int <= to_signed(-798,32);
				when 1626 => sin_data_int <= to_signed(603,32); cos_data_int <= to_signed(-799,32);
				when 1627 => sin_data_int <= to_signed(602,32); cos_data_int <= to_signed(-800,32);
				when 1628 => sin_data_int <= to_signed(601,32); cos_data_int <= to_signed(-800,32);
				when 1629 => sin_data_int <= to_signed(599,32); cos_data_int <= to_signed(-801,32);
				when 1630 => sin_data_int <= to_signed(598,32); cos_data_int <= to_signed(-802,32);
				when 1631 => sin_data_int <= to_signed(597,32); cos_data_int <= to_signed(-803,32);
				when 1632 => sin_data_int <= to_signed(596,32); cos_data_int <= to_signed(-804,32);
				when 1633 => sin_data_int <= to_signed(594,32); cos_data_int <= to_signed(-805,32);
				when 1634 => sin_data_int <= to_signed(593,32); cos_data_int <= to_signed(-806,32);
				when 1635 => sin_data_int <= to_signed(592,32); cos_data_int <= to_signed(-807,32);
				when 1636 => sin_data_int <= to_signed(591,32); cos_data_int <= to_signed(-808,32);
				when 1637 => sin_data_int <= to_signed(590,32); cos_data_int <= to_signed(-809,32);
				when 1638 => sin_data_int <= to_signed(588,32); cos_data_int <= to_signed(-810,32);
				when 1639 => sin_data_int <= to_signed(587,32); cos_data_int <= to_signed(-810,32);
				when 1640 => sin_data_int <= to_signed(586,32); cos_data_int <= to_signed(-811,32);
				when 1641 => sin_data_int <= to_signed(585,32); cos_data_int <= to_signed(-812,32);
				when 1642 => sin_data_int <= to_signed(583,32); cos_data_int <= to_signed(-813,32);
				when 1643 => sin_data_int <= to_signed(582,32); cos_data_int <= to_signed(-814,32);
				when 1644 => sin_data_int <= to_signed(581,32); cos_data_int <= to_signed(-815,32);
				when 1645 => sin_data_int <= to_signed(580,32); cos_data_int <= to_signed(-816,32);
				when 1646 => sin_data_int <= to_signed(578,32); cos_data_int <= to_signed(-817,32);
				when 1647 => sin_data_int <= to_signed(577,32); cos_data_int <= to_signed(-818,32);
				when 1648 => sin_data_int <= to_signed(576,32); cos_data_int <= to_signed(-818,32);
				when 1649 => sin_data_int <= to_signed(575,32); cos_data_int <= to_signed(-819,32);
				when 1650 => sin_data_int <= to_signed(573,32); cos_data_int <= to_signed(-820,32);
				when 1651 => sin_data_int <= to_signed(572,32); cos_data_int <= to_signed(-821,32);
				when 1652 => sin_data_int <= to_signed(571,32); cos_data_int <= to_signed(-822,32);
				when 1653 => sin_data_int <= to_signed(570,32); cos_data_int <= to_signed(-823,32);
				when 1654 => sin_data_int <= to_signed(568,32); cos_data_int <= to_signed(-824,32);
				when 1655 => sin_data_int <= to_signed(567,32); cos_data_int <= to_signed(-825,32);
				when 1656 => sin_data_int <= to_signed(566,32); cos_data_int <= to_signed(-825,32);
				when 1657 => sin_data_int <= to_signed(564,32); cos_data_int <= to_signed(-826,32);
				when 1658 => sin_data_int <= to_signed(563,32); cos_data_int <= to_signed(-827,32);
				when 1659 => sin_data_int <= to_signed(562,32); cos_data_int <= to_signed(-828,32);
				when 1660 => sin_data_int <= to_signed(561,32); cos_data_int <= to_signed(-829,32);
				when 1661 => sin_data_int <= to_signed(559,32); cos_data_int <= to_signed(-830,32);
				when 1662 => sin_data_int <= to_signed(558,32); cos_data_int <= to_signed(-831,32);
				when 1663 => sin_data_int <= to_signed(557,32); cos_data_int <= to_signed(-831,32);
				when 1664 => sin_data_int <= to_signed(556,32); cos_data_int <= to_signed(-832,32);
				when 1665 => sin_data_int <= to_signed(554,32); cos_data_int <= to_signed(-833,32);
				when 1666 => sin_data_int <= to_signed(553,32); cos_data_int <= to_signed(-834,32);
				when 1667 => sin_data_int <= to_signed(552,32); cos_data_int <= to_signed(-835,32);
				when 1668 => sin_data_int <= to_signed(550,32); cos_data_int <= to_signed(-836,32);
				when 1669 => sin_data_int <= to_signed(549,32); cos_data_int <= to_signed(-837,32);
				when 1670 => sin_data_int <= to_signed(548,32); cos_data_int <= to_signed(-837,32);
				when 1671 => sin_data_int <= to_signed(547,32); cos_data_int <= to_signed(-838,32);
				when 1672 => sin_data_int <= to_signed(545,32); cos_data_int <= to_signed(-839,32);
				when 1673 => sin_data_int <= to_signed(544,32); cos_data_int <= to_signed(-840,32);
				when 1674 => sin_data_int <= to_signed(543,32); cos_data_int <= to_signed(-841,32);
				when 1675 => sin_data_int <= to_signed(541,32); cos_data_int <= to_signed(-842,32);
				when 1676 => sin_data_int <= to_signed(540,32); cos_data_int <= to_signed(-842,32);
				when 1677 => sin_data_int <= to_signed(539,32); cos_data_int <= to_signed(-843,32);
				when 1678 => sin_data_int <= to_signed(538,32); cos_data_int <= to_signed(-844,32);
				when 1679 => sin_data_int <= to_signed(536,32); cos_data_int <= to_signed(-845,32);
				when 1680 => sin_data_int <= to_signed(535,32); cos_data_int <= to_signed(-846,32);
				when 1681 => sin_data_int <= to_signed(534,32); cos_data_int <= to_signed(-846,32);
				when 1682 => sin_data_int <= to_signed(532,32); cos_data_int <= to_signed(-847,32);
				when 1683 => sin_data_int <= to_signed(531,32); cos_data_int <= to_signed(-848,32);
				when 1684 => sin_data_int <= to_signed(530,32); cos_data_int <= to_signed(-849,32);
				when 1685 => sin_data_int <= to_signed(529,32); cos_data_int <= to_signed(-850,32);
				when 1686 => sin_data_int <= to_signed(527,32); cos_data_int <= to_signed(-851,32);
				when 1687 => sin_data_int <= to_signed(526,32); cos_data_int <= to_signed(-851,32);
				when 1688 => sin_data_int <= to_signed(525,32); cos_data_int <= to_signed(-852,32);
				when 1689 => sin_data_int <= to_signed(523,32); cos_data_int <= to_signed(-853,32);
				when 1690 => sin_data_int <= to_signed(522,32); cos_data_int <= to_signed(-854,32);
				when 1691 => sin_data_int <= to_signed(521,32); cos_data_int <= to_signed(-855,32);
				when 1692 => sin_data_int <= to_signed(519,32); cos_data_int <= to_signed(-855,32);
				when 1693 => sin_data_int <= to_signed(518,32); cos_data_int <= to_signed(-856,32);
				when 1694 => sin_data_int <= to_signed(517,32); cos_data_int <= to_signed(-857,32);
				when 1695 => sin_data_int <= to_signed(515,32); cos_data_int <= to_signed(-858,32);
				when 1696 => sin_data_int <= to_signed(514,32); cos_data_int <= to_signed(-859,32);
				when 1697 => sin_data_int <= to_signed(513,32); cos_data_int <= to_signed(-859,32);
				when 1698 => sin_data_int <= to_signed(511,32); cos_data_int <= to_signed(-860,32);
				when 1699 => sin_data_int <= to_signed(510,32); cos_data_int <= to_signed(-861,32);
				when 1700 => sin_data_int <= to_signed(509,32); cos_data_int <= to_signed(-862,32);
				when 1701 => sin_data_int <= to_signed(508,32); cos_data_int <= to_signed(-862,32);
				when 1702 => sin_data_int <= to_signed(506,32); cos_data_int <= to_signed(-863,32);
				when 1703 => sin_data_int <= to_signed(505,32); cos_data_int <= to_signed(-864,32);
				when 1704 => sin_data_int <= to_signed(504,32); cos_data_int <= to_signed(-865,32);
				when 1705 => sin_data_int <= to_signed(502,32); cos_data_int <= to_signed(-866,32);
				when 1706 => sin_data_int <= to_signed(501,32); cos_data_int <= to_signed(-866,32);
				when 1707 => sin_data_int <= to_signed(500,32); cos_data_int <= to_signed(-867,32);
				when 1708 => sin_data_int <= to_signed(498,32); cos_data_int <= to_signed(-868,32);
				when 1709 => sin_data_int <= to_signed(497,32); cos_data_int <= to_signed(-869,32);
				when 1710 => sin_data_int <= to_signed(496,32); cos_data_int <= to_signed(-869,32);
				when 1711 => sin_data_int <= to_signed(494,32); cos_data_int <= to_signed(-870,32);
				when 1712 => sin_data_int <= to_signed(493,32); cos_data_int <= to_signed(-871,32);
				when 1713 => sin_data_int <= to_signed(492,32); cos_data_int <= to_signed(-872,32);
				when 1714 => sin_data_int <= to_signed(490,32); cos_data_int <= to_signed(-872,32);
				when 1715 => sin_data_int <= to_signed(489,32); cos_data_int <= to_signed(-873,32);
				when 1716 => sin_data_int <= to_signed(488,32); cos_data_int <= to_signed(-874,32);
				when 1717 => sin_data_int <= to_signed(486,32); cos_data_int <= to_signed(-875,32);
				when 1718 => sin_data_int <= to_signed(485,32); cos_data_int <= to_signed(-875,32);
				when 1719 => sin_data_int <= to_signed(484,32); cos_data_int <= to_signed(-876,32);
				when 1720 => sin_data_int <= to_signed(482,32); cos_data_int <= to_signed(-877,32);
				when 1721 => sin_data_int <= to_signed(481,32); cos_data_int <= to_signed(-878,32);
				when 1722 => sin_data_int <= to_signed(479,32); cos_data_int <= to_signed(-878,32);
				when 1723 => sin_data_int <= to_signed(478,32); cos_data_int <= to_signed(-879,32);
				when 1724 => sin_data_int <= to_signed(477,32); cos_data_int <= to_signed(-880,32);
				when 1725 => sin_data_int <= to_signed(475,32); cos_data_int <= to_signed(-880,32);
				when 1726 => sin_data_int <= to_signed(474,32); cos_data_int <= to_signed(-881,32);
				when 1727 => sin_data_int <= to_signed(473,32); cos_data_int <= to_signed(-882,32);
				when 1728 => sin_data_int <= to_signed(471,32); cos_data_int <= to_signed(-883,32);
				when 1729 => sin_data_int <= to_signed(470,32); cos_data_int <= to_signed(-883,32);
				when 1730 => sin_data_int <= to_signed(469,32); cos_data_int <= to_signed(-884,32);
				when 1731 => sin_data_int <= to_signed(467,32); cos_data_int <= to_signed(-885,32);
				when 1732 => sin_data_int <= to_signed(466,32); cos_data_int <= to_signed(-886,32);
				when 1733 => sin_data_int <= to_signed(465,32); cos_data_int <= to_signed(-886,32);
				when 1734 => sin_data_int <= to_signed(463,32); cos_data_int <= to_signed(-887,32);
				when 1735 => sin_data_int <= to_signed(462,32); cos_data_int <= to_signed(-888,32);
				when 1736 => sin_data_int <= to_signed(461,32); cos_data_int <= to_signed(-888,32);
				when 1737 => sin_data_int <= to_signed(459,32); cos_data_int <= to_signed(-889,32);
				when 1738 => sin_data_int <= to_signed(458,32); cos_data_int <= to_signed(-890,32);
				when 1739 => sin_data_int <= to_signed(456,32); cos_data_int <= to_signed(-890,32);
				when 1740 => sin_data_int <= to_signed(455,32); cos_data_int <= to_signed(-891,32);
				when 1741 => sin_data_int <= to_signed(454,32); cos_data_int <= to_signed(-892,32);
				when 1742 => sin_data_int <= to_signed(452,32); cos_data_int <= to_signed(-893,32);
				when 1743 => sin_data_int <= to_signed(451,32); cos_data_int <= to_signed(-893,32);
				when 1744 => sin_data_int <= to_signed(450,32); cos_data_int <= to_signed(-894,32);
				when 1745 => sin_data_int <= to_signed(448,32); cos_data_int <= to_signed(-895,32);
				when 1746 => sin_data_int <= to_signed(447,32); cos_data_int <= to_signed(-895,32);
				when 1747 => sin_data_int <= to_signed(445,32); cos_data_int <= to_signed(-896,32);
				when 1748 => sin_data_int <= to_signed(444,32); cos_data_int <= to_signed(-897,32);
				when 1749 => sin_data_int <= to_signed(443,32); cos_data_int <= to_signed(-897,32);
				when 1750 => sin_data_int <= to_signed(441,32); cos_data_int <= to_signed(-898,32);
				when 1751 => sin_data_int <= to_signed(440,32); cos_data_int <= to_signed(-899,32);
				when 1752 => sin_data_int <= to_signed(439,32); cos_data_int <= to_signed(-899,32);
				when 1753 => sin_data_int <= to_signed(437,32); cos_data_int <= to_signed(-900,32);
				when 1754 => sin_data_int <= to_signed(436,32); cos_data_int <= to_signed(-901,32);
				when 1755 => sin_data_int <= to_signed(434,32); cos_data_int <= to_signed(-901,32);
				when 1756 => sin_data_int <= to_signed(433,32); cos_data_int <= to_signed(-902,32);
				when 1757 => sin_data_int <= to_signed(432,32); cos_data_int <= to_signed(-903,32);
				when 1758 => sin_data_int <= to_signed(430,32); cos_data_int <= to_signed(-903,32);
				when 1759 => sin_data_int <= to_signed(429,32); cos_data_int <= to_signed(-904,32);
				when 1760 => sin_data_int <= to_signed(428,32); cos_data_int <= to_signed(-905,32);
				when 1761 => sin_data_int <= to_signed(426,32); cos_data_int <= to_signed(-905,32);
				when 1762 => sin_data_int <= to_signed(425,32); cos_data_int <= to_signed(-906,32);
				when 1763 => sin_data_int <= to_signed(423,32); cos_data_int <= to_signed(-907,32);
				when 1764 => sin_data_int <= to_signed(422,32); cos_data_int <= to_signed(-907,32);
				when 1765 => sin_data_int <= to_signed(421,32); cos_data_int <= to_signed(-908,32);
				when 1766 => sin_data_int <= to_signed(419,32); cos_data_int <= to_signed(-909,32);
				when 1767 => sin_data_int <= to_signed(418,32); cos_data_int <= to_signed(-909,32);
				when 1768 => sin_data_int <= to_signed(416,32); cos_data_int <= to_signed(-910,32);
				when 1769 => sin_data_int <= to_signed(415,32); cos_data_int <= to_signed(-910,32);
				when 1770 => sin_data_int <= to_signed(414,32); cos_data_int <= to_signed(-911,32);
				when 1771 => sin_data_int <= to_signed(412,32); cos_data_int <= to_signed(-912,32);
				when 1772 => sin_data_int <= to_signed(411,32); cos_data_int <= to_signed(-912,32);
				when 1773 => sin_data_int <= to_signed(409,32); cos_data_int <= to_signed(-913,32);
				when 1774 => sin_data_int <= to_signed(408,32); cos_data_int <= to_signed(-914,32);
				when 1775 => sin_data_int <= to_signed(407,32); cos_data_int <= to_signed(-914,32);
				when 1776 => sin_data_int <= to_signed(405,32); cos_data_int <= to_signed(-915,32);
				when 1777 => sin_data_int <= to_signed(404,32); cos_data_int <= to_signed(-915,32);
				when 1778 => sin_data_int <= to_signed(402,32); cos_data_int <= to_signed(-916,32);
				when 1779 => sin_data_int <= to_signed(401,32); cos_data_int <= to_signed(-917,32);
				when 1780 => sin_data_int <= to_signed(400,32); cos_data_int <= to_signed(-917,32);
				when 1781 => sin_data_int <= to_signed(398,32); cos_data_int <= to_signed(-918,32);
				when 1782 => sin_data_int <= to_signed(397,32); cos_data_int <= to_signed(-919,32);
				when 1783 => sin_data_int <= to_signed(395,32); cos_data_int <= to_signed(-919,32);
				when 1784 => sin_data_int <= to_signed(394,32); cos_data_int <= to_signed(-920,32);
				when 1785 => sin_data_int <= to_signed(393,32); cos_data_int <= to_signed(-920,32);
				when 1786 => sin_data_int <= to_signed(391,32); cos_data_int <= to_signed(-921,32);
				when 1787 => sin_data_int <= to_signed(390,32); cos_data_int <= to_signed(-922,32);
				when 1788 => sin_data_int <= to_signed(388,32); cos_data_int <= to_signed(-922,32);
				when 1789 => sin_data_int <= to_signed(387,32); cos_data_int <= to_signed(-923,32);
				when 1790 => sin_data_int <= to_signed(386,32); cos_data_int <= to_signed(-923,32);
				when 1791 => sin_data_int <= to_signed(384,32); cos_data_int <= to_signed(-924,32);
				when 1792 => sin_data_int <= to_signed(383,32); cos_data_int <= to_signed(-924,32);
				when 1793 => sin_data_int <= to_signed(381,32); cos_data_int <= to_signed(-925,32);
				when 1794 => sin_data_int <= to_signed(380,32); cos_data_int <= to_signed(-926,32);
				when 1795 => sin_data_int <= to_signed(378,32); cos_data_int <= to_signed(-926,32);
				when 1796 => sin_data_int <= to_signed(377,32); cos_data_int <= to_signed(-927,32);
				when 1797 => sin_data_int <= to_signed(376,32); cos_data_int <= to_signed(-927,32);
				when 1798 => sin_data_int <= to_signed(374,32); cos_data_int <= to_signed(-928,32);
				when 1799 => sin_data_int <= to_signed(373,32); cos_data_int <= to_signed(-929,32);
				when 1800 => sin_data_int <= to_signed(371,32); cos_data_int <= to_signed(-929,32);
				when 1801 => sin_data_int <= to_signed(370,32); cos_data_int <= to_signed(-930,32);
				when 1802 => sin_data_int <= to_signed(368,32); cos_data_int <= to_signed(-930,32);
				when 1803 => sin_data_int <= to_signed(367,32); cos_data_int <= to_signed(-931,32);
				when 1804 => sin_data_int <= to_signed(366,32); cos_data_int <= to_signed(-931,32);
				when 1805 => sin_data_int <= to_signed(364,32); cos_data_int <= to_signed(-932,32);
				when 1806 => sin_data_int <= to_signed(363,32); cos_data_int <= to_signed(-932,32);
				when 1807 => sin_data_int <= to_signed(361,32); cos_data_int <= to_signed(-933,32);
				when 1808 => sin_data_int <= to_signed(360,32); cos_data_int <= to_signed(-934,32);
				when 1809 => sin_data_int <= to_signed(358,32); cos_data_int <= to_signed(-934,32);
				when 1810 => sin_data_int <= to_signed(357,32); cos_data_int <= to_signed(-935,32);
				when 1811 => sin_data_int <= to_signed(356,32); cos_data_int <= to_signed(-935,32);
				when 1812 => sin_data_int <= to_signed(354,32); cos_data_int <= to_signed(-936,32);
				when 1813 => sin_data_int <= to_signed(353,32); cos_data_int <= to_signed(-936,32);
				when 1814 => sin_data_int <= to_signed(351,32); cos_data_int <= to_signed(-937,32);
				when 1815 => sin_data_int <= to_signed(350,32); cos_data_int <= to_signed(-937,32);
				when 1816 => sin_data_int <= to_signed(348,32); cos_data_int <= to_signed(-938,32);
				when 1817 => sin_data_int <= to_signed(347,32); cos_data_int <= to_signed(-938,32);
				when 1818 => sin_data_int <= to_signed(346,32); cos_data_int <= to_signed(-939,32);
				when 1819 => sin_data_int <= to_signed(344,32); cos_data_int <= to_signed(-939,32);
				when 1820 => sin_data_int <= to_signed(343,32); cos_data_int <= to_signed(-940,32);
				when 1821 => sin_data_int <= to_signed(341,32); cos_data_int <= to_signed(-941,32);
				when 1822 => sin_data_int <= to_signed(340,32); cos_data_int <= to_signed(-941,32);
				when 1823 => sin_data_int <= to_signed(338,32); cos_data_int <= to_signed(-942,32);
				when 1824 => sin_data_int <= to_signed(337,32); cos_data_int <= to_signed(-942,32);
				when 1825 => sin_data_int <= to_signed(335,32); cos_data_int <= to_signed(-943,32);
				when 1826 => sin_data_int <= to_signed(334,32); cos_data_int <= to_signed(-943,32);
				when 1827 => sin_data_int <= to_signed(333,32); cos_data_int <= to_signed(-944,32);
				when 1828 => sin_data_int <= to_signed(331,32); cos_data_int <= to_signed(-944,32);
				when 1829 => sin_data_int <= to_signed(330,32); cos_data_int <= to_signed(-945,32);
				when 1830 => sin_data_int <= to_signed(328,32); cos_data_int <= to_signed(-945,32);
				when 1831 => sin_data_int <= to_signed(327,32); cos_data_int <= to_signed(-946,32);
				when 1832 => sin_data_int <= to_signed(325,32); cos_data_int <= to_signed(-946,32);
				when 1833 => sin_data_int <= to_signed(324,32); cos_data_int <= to_signed(-947,32);
				when 1834 => sin_data_int <= to_signed(322,32); cos_data_int <= to_signed(-947,32);
				when 1835 => sin_data_int <= to_signed(321,32); cos_data_int <= to_signed(-948,32);
				when 1836 => sin_data_int <= to_signed(320,32); cos_data_int <= to_signed(-948,32);
				when 1837 => sin_data_int <= to_signed(318,32); cos_data_int <= to_signed(-949,32);
				when 1838 => sin_data_int <= to_signed(317,32); cos_data_int <= to_signed(-949,32);
				when 1839 => sin_data_int <= to_signed(315,32); cos_data_int <= to_signed(-950,32);
				when 1840 => sin_data_int <= to_signed(314,32); cos_data_int <= to_signed(-950,32);
				when 1841 => sin_data_int <= to_signed(312,32); cos_data_int <= to_signed(-950,32);
				when 1842 => sin_data_int <= to_signed(311,32); cos_data_int <= to_signed(-951,32);
				when 1843 => sin_data_int <= to_signed(309,32); cos_data_int <= to_signed(-951,32);
				when 1844 => sin_data_int <= to_signed(308,32); cos_data_int <= to_signed(-952,32);
				when 1845 => sin_data_int <= to_signed(306,32); cos_data_int <= to_signed(-952,32);
				when 1846 => sin_data_int <= to_signed(305,32); cos_data_int <= to_signed(-953,32);
				when 1847 => sin_data_int <= to_signed(303,32); cos_data_int <= to_signed(-953,32);
				when 1848 => sin_data_int <= to_signed(302,32); cos_data_int <= to_signed(-954,32);
				when 1849 => sin_data_int <= to_signed(301,32); cos_data_int <= to_signed(-954,32);
				when 1850 => sin_data_int <= to_signed(299,32); cos_data_int <= to_signed(-955,32);
				when 1851 => sin_data_int <= to_signed(298,32); cos_data_int <= to_signed(-955,32);
				when 1852 => sin_data_int <= to_signed(296,32); cos_data_int <= to_signed(-956,32);
				when 1853 => sin_data_int <= to_signed(295,32); cos_data_int <= to_signed(-956,32);
				when 1854 => sin_data_int <= to_signed(293,32); cos_data_int <= to_signed(-956,32);
				when 1855 => sin_data_int <= to_signed(292,32); cos_data_int <= to_signed(-957,32);
				when 1856 => sin_data_int <= to_signed(290,32); cos_data_int <= to_signed(-957,32);
				when 1857 => sin_data_int <= to_signed(289,32); cos_data_int <= to_signed(-958,32);
				when 1858 => sin_data_int <= to_signed(287,32); cos_data_int <= to_signed(-958,32);
				when 1859 => sin_data_int <= to_signed(286,32); cos_data_int <= to_signed(-959,32);
				when 1860 => sin_data_int <= to_signed(284,32); cos_data_int <= to_signed(-959,32);
				when 1861 => sin_data_int <= to_signed(283,32); cos_data_int <= to_signed(-960,32);
				when 1862 => sin_data_int <= to_signed(281,32); cos_data_int <= to_signed(-960,32);
				when 1863 => sin_data_int <= to_signed(280,32); cos_data_int <= to_signed(-960,32);
				when 1864 => sin_data_int <= to_signed(279,32); cos_data_int <= to_signed(-961,32);
				when 1865 => sin_data_int <= to_signed(277,32); cos_data_int <= to_signed(-961,32);
				when 1866 => sin_data_int <= to_signed(276,32); cos_data_int <= to_signed(-962,32);
				when 1867 => sin_data_int <= to_signed(274,32); cos_data_int <= to_signed(-962,32);
				when 1868 => sin_data_int <= to_signed(273,32); cos_data_int <= to_signed(-963,32);
				when 1869 => sin_data_int <= to_signed(271,32); cos_data_int <= to_signed(-963,32);
				when 1870 => sin_data_int <= to_signed(270,32); cos_data_int <= to_signed(-963,32);
				when 1871 => sin_data_int <= to_signed(268,32); cos_data_int <= to_signed(-964,32);
				when 1872 => sin_data_int <= to_signed(267,32); cos_data_int <= to_signed(-964,32);
				when 1873 => sin_data_int <= to_signed(265,32); cos_data_int <= to_signed(-965,32);
				when 1874 => sin_data_int <= to_signed(264,32); cos_data_int <= to_signed(-965,32);
				when 1875 => sin_data_int <= to_signed(262,32); cos_data_int <= to_signed(-965,32);
				when 1876 => sin_data_int <= to_signed(261,32); cos_data_int <= to_signed(-966,32);
				when 1877 => sin_data_int <= to_signed(259,32); cos_data_int <= to_signed(-966,32);
				when 1878 => sin_data_int <= to_signed(258,32); cos_data_int <= to_signed(-967,32);
				when 1879 => sin_data_int <= to_signed(256,32); cos_data_int <= to_signed(-967,32);
				when 1880 => sin_data_int <= to_signed(255,32); cos_data_int <= to_signed(-967,32);
				when 1881 => sin_data_int <= to_signed(253,32); cos_data_int <= to_signed(-968,32);
				when 1882 => sin_data_int <= to_signed(252,32); cos_data_int <= to_signed(-968,32);
				when 1883 => sin_data_int <= to_signed(250,32); cos_data_int <= to_signed(-969,32);
				when 1884 => sin_data_int <= to_signed(249,32); cos_data_int <= to_signed(-969,32);
				when 1885 => sin_data_int <= to_signed(247,32); cos_data_int <= to_signed(-969,32);
				when 1886 => sin_data_int <= to_signed(246,32); cos_data_int <= to_signed(-970,32);
				when 1887 => sin_data_int <= to_signed(244,32); cos_data_int <= to_signed(-970,32);
				when 1888 => sin_data_int <= to_signed(243,32); cos_data_int <= to_signed(-970,32);
				when 1889 => sin_data_int <= to_signed(241,32); cos_data_int <= to_signed(-971,32);
				when 1890 => sin_data_int <= to_signed(240,32); cos_data_int <= to_signed(-971,32);
				when 1891 => sin_data_int <= to_signed(239,32); cos_data_int <= to_signed(-972,32);
				when 1892 => sin_data_int <= to_signed(237,32); cos_data_int <= to_signed(-972,32);
				when 1893 => sin_data_int <= to_signed(236,32); cos_data_int <= to_signed(-972,32);
				when 1894 => sin_data_int <= to_signed(234,32); cos_data_int <= to_signed(-973,32);
				when 1895 => sin_data_int <= to_signed(233,32); cos_data_int <= to_signed(-973,32);
				when 1896 => sin_data_int <= to_signed(231,32); cos_data_int <= to_signed(-973,32);
				when 1897 => sin_data_int <= to_signed(230,32); cos_data_int <= to_signed(-974,32);
				when 1898 => sin_data_int <= to_signed(228,32); cos_data_int <= to_signed(-974,32);
				when 1899 => sin_data_int <= to_signed(227,32); cos_data_int <= to_signed(-974,32);
				when 1900 => sin_data_int <= to_signed(225,32); cos_data_int <= to_signed(-975,32);
				when 1901 => sin_data_int <= to_signed(224,32); cos_data_int <= to_signed(-975,32);
				when 1902 => sin_data_int <= to_signed(222,32); cos_data_int <= to_signed(-975,32);
				when 1903 => sin_data_int <= to_signed(221,32); cos_data_int <= to_signed(-976,32);
				when 1904 => sin_data_int <= to_signed(219,32); cos_data_int <= to_signed(-976,32);
				when 1905 => sin_data_int <= to_signed(218,32); cos_data_int <= to_signed(-976,32);
				when 1906 => sin_data_int <= to_signed(216,32); cos_data_int <= to_signed(-977,32);
				when 1907 => sin_data_int <= to_signed(215,32); cos_data_int <= to_signed(-977,32);
				when 1908 => sin_data_int <= to_signed(213,32); cos_data_int <= to_signed(-977,32);
				when 1909 => sin_data_int <= to_signed(212,32); cos_data_int <= to_signed(-978,32);
				when 1910 => sin_data_int <= to_signed(210,32); cos_data_int <= to_signed(-978,32);
				when 1911 => sin_data_int <= to_signed(209,32); cos_data_int <= to_signed(-978,32);
				when 1912 => sin_data_int <= to_signed(207,32); cos_data_int <= to_signed(-979,32);
				when 1913 => sin_data_int <= to_signed(206,32); cos_data_int <= to_signed(-979,32);
				when 1914 => sin_data_int <= to_signed(204,32); cos_data_int <= to_signed(-979,32);
				when 1915 => sin_data_int <= to_signed(203,32); cos_data_int <= to_signed(-980,32);
				when 1916 => sin_data_int <= to_signed(201,32); cos_data_int <= to_signed(-980,32);
				when 1917 => sin_data_int <= to_signed(200,32); cos_data_int <= to_signed(-980,32);
				when 1918 => sin_data_int <= to_signed(198,32); cos_data_int <= to_signed(-980,32);
				when 1919 => sin_data_int <= to_signed(197,32); cos_data_int <= to_signed(-981,32);
				when 1920 => sin_data_int <= to_signed(195,32); cos_data_int <= to_signed(-981,32);
				when 1921 => sin_data_int <= to_signed(194,32); cos_data_int <= to_signed(-981,32);
				when 1922 => sin_data_int <= to_signed(192,32); cos_data_int <= to_signed(-982,32);
				when 1923 => sin_data_int <= to_signed(191,32); cos_data_int <= to_signed(-982,32);
				when 1924 => sin_data_int <= to_signed(189,32); cos_data_int <= to_signed(-982,32);
				when 1925 => sin_data_int <= to_signed(188,32); cos_data_int <= to_signed(-983,32);
				when 1926 => sin_data_int <= to_signed(186,32); cos_data_int <= to_signed(-983,32);
				when 1927 => sin_data_int <= to_signed(185,32); cos_data_int <= to_signed(-983,32);
				when 1928 => sin_data_int <= to_signed(183,32); cos_data_int <= to_signed(-983,32);
				when 1929 => sin_data_int <= to_signed(182,32); cos_data_int <= to_signed(-984,32);
				when 1930 => sin_data_int <= to_signed(180,32); cos_data_int <= to_signed(-984,32);
				when 1931 => sin_data_int <= to_signed(179,32); cos_data_int <= to_signed(-984,32);
				when 1932 => sin_data_int <= to_signed(177,32); cos_data_int <= to_signed(-984,32);
				when 1933 => sin_data_int <= to_signed(175,32); cos_data_int <= to_signed(-985,32);
				when 1934 => sin_data_int <= to_signed(174,32); cos_data_int <= to_signed(-985,32);
				when 1935 => sin_data_int <= to_signed(172,32); cos_data_int <= to_signed(-985,32);
				when 1936 => sin_data_int <= to_signed(171,32); cos_data_int <= to_signed(-986,32);
				when 1937 => sin_data_int <= to_signed(169,32); cos_data_int <= to_signed(-986,32);
				when 1938 => sin_data_int <= to_signed(168,32); cos_data_int <= to_signed(-986,32);
				when 1939 => sin_data_int <= to_signed(166,32); cos_data_int <= to_signed(-986,32);
				when 1940 => sin_data_int <= to_signed(165,32); cos_data_int <= to_signed(-987,32);
				when 1941 => sin_data_int <= to_signed(163,32); cos_data_int <= to_signed(-987,32);
				when 1942 => sin_data_int <= to_signed(162,32); cos_data_int <= to_signed(-987,32);
				when 1943 => sin_data_int <= to_signed(160,32); cos_data_int <= to_signed(-987,32);
				when 1944 => sin_data_int <= to_signed(159,32); cos_data_int <= to_signed(-988,32);
				when 1945 => sin_data_int <= to_signed(157,32); cos_data_int <= to_signed(-988,32);
				when 1946 => sin_data_int <= to_signed(156,32); cos_data_int <= to_signed(-988,32);
				when 1947 => sin_data_int <= to_signed(154,32); cos_data_int <= to_signed(-988,32);
				when 1948 => sin_data_int <= to_signed(153,32); cos_data_int <= to_signed(-988,32);
				when 1949 => sin_data_int <= to_signed(151,32); cos_data_int <= to_signed(-989,32);
				when 1950 => sin_data_int <= to_signed(150,32); cos_data_int <= to_signed(-989,32);
				when 1951 => sin_data_int <= to_signed(148,32); cos_data_int <= to_signed(-989,32);
				when 1952 => sin_data_int <= to_signed(147,32); cos_data_int <= to_signed(-989,32);
				when 1953 => sin_data_int <= to_signed(145,32); cos_data_int <= to_signed(-990,32);
				when 1954 => sin_data_int <= to_signed(144,32); cos_data_int <= to_signed(-990,32);
				when 1955 => sin_data_int <= to_signed(142,32); cos_data_int <= to_signed(-990,32);
				when 1956 => sin_data_int <= to_signed(141,32); cos_data_int <= to_signed(-990,32);
				when 1957 => sin_data_int <= to_signed(139,32); cos_data_int <= to_signed(-990,32);
				when 1958 => sin_data_int <= to_signed(138,32); cos_data_int <= to_signed(-991,32);
				when 1959 => sin_data_int <= to_signed(136,32); cos_data_int <= to_signed(-991,32);
				when 1960 => sin_data_int <= to_signed(135,32); cos_data_int <= to_signed(-991,32);
				when 1961 => sin_data_int <= to_signed(133,32); cos_data_int <= to_signed(-991,32);
				when 1962 => sin_data_int <= to_signed(132,32); cos_data_int <= to_signed(-992,32);
				when 1963 => sin_data_int <= to_signed(130,32); cos_data_int <= to_signed(-992,32);
				when 1964 => sin_data_int <= to_signed(128,32); cos_data_int <= to_signed(-992,32);
				when 1965 => sin_data_int <= to_signed(127,32); cos_data_int <= to_signed(-992,32);
				when 1966 => sin_data_int <= to_signed(125,32); cos_data_int <= to_signed(-992,32);
				when 1967 => sin_data_int <= to_signed(124,32); cos_data_int <= to_signed(-992,32);
				when 1968 => sin_data_int <= to_signed(122,32); cos_data_int <= to_signed(-993,32);
				when 1969 => sin_data_int <= to_signed(121,32); cos_data_int <= to_signed(-993,32);
				when 1970 => sin_data_int <= to_signed(119,32); cos_data_int <= to_signed(-993,32);
				when 1971 => sin_data_int <= to_signed(118,32); cos_data_int <= to_signed(-993,32);
				when 1972 => sin_data_int <= to_signed(116,32); cos_data_int <= to_signed(-993,32);
				when 1973 => sin_data_int <= to_signed(115,32); cos_data_int <= to_signed(-994,32);
				when 1974 => sin_data_int <= to_signed(113,32); cos_data_int <= to_signed(-994,32);
				when 1975 => sin_data_int <= to_signed(112,32); cos_data_int <= to_signed(-994,32);
				when 1976 => sin_data_int <= to_signed(110,32); cos_data_int <= to_signed(-994,32);
				when 1977 => sin_data_int <= to_signed(109,32); cos_data_int <= to_signed(-994,32);
				when 1978 => sin_data_int <= to_signed(107,32); cos_data_int <= to_signed(-994,32);
				when 1979 => sin_data_int <= to_signed(106,32); cos_data_int <= to_signed(-995,32);
				when 1980 => sin_data_int <= to_signed(104,32); cos_data_int <= to_signed(-995,32);
				when 1981 => sin_data_int <= to_signed(103,32); cos_data_int <= to_signed(-995,32);
				when 1982 => sin_data_int <= to_signed(101,32); cos_data_int <= to_signed(-995,32);
				when 1983 => sin_data_int <= to_signed(100,32); cos_data_int <= to_signed(-995,32);
				when 1984 => sin_data_int <= to_signed(98,32); cos_data_int <= to_signed(-995,32);
				when 1985 => sin_data_int <= to_signed(96,32); cos_data_int <= to_signed(-995,32);
				when 1986 => sin_data_int <= to_signed(95,32); cos_data_int <= to_signed(-996,32);
				when 1987 => sin_data_int <= to_signed(93,32); cos_data_int <= to_signed(-996,32);
				when 1988 => sin_data_int <= to_signed(92,32); cos_data_int <= to_signed(-996,32);
				when 1989 => sin_data_int <= to_signed(90,32); cos_data_int <= to_signed(-996,32);
				when 1990 => sin_data_int <= to_signed(89,32); cos_data_int <= to_signed(-996,32);
				when 1991 => sin_data_int <= to_signed(87,32); cos_data_int <= to_signed(-996,32);
				when 1992 => sin_data_int <= to_signed(86,32); cos_data_int <= to_signed(-996,32);
				when 1993 => sin_data_int <= to_signed(84,32); cos_data_int <= to_signed(-997,32);
				when 1994 => sin_data_int <= to_signed(83,32); cos_data_int <= to_signed(-997,32);
				when 1995 => sin_data_int <= to_signed(81,32); cos_data_int <= to_signed(-997,32);
				when 1996 => sin_data_int <= to_signed(80,32); cos_data_int <= to_signed(-997,32);
				when 1997 => sin_data_int <= to_signed(78,32); cos_data_int <= to_signed(-997,32);
				when 1998 => sin_data_int <= to_signed(77,32); cos_data_int <= to_signed(-997,32);
				when 1999 => sin_data_int <= to_signed(75,32); cos_data_int <= to_signed(-997,32);
				when 2000 => sin_data_int <= to_signed(74,32); cos_data_int <= to_signed(-997,32);
				when 2001 => sin_data_int <= to_signed(72,32); cos_data_int <= to_signed(-998,32);
				when 2002 => sin_data_int <= to_signed(71,32); cos_data_int <= to_signed(-998,32);
				when 2003 => sin_data_int <= to_signed(69,32); cos_data_int <= to_signed(-998,32);
				when 2004 => sin_data_int <= to_signed(67,32); cos_data_int <= to_signed(-998,32);
				when 2005 => sin_data_int <= to_signed(66,32); cos_data_int <= to_signed(-998,32);
				when 2006 => sin_data_int <= to_signed(64,32); cos_data_int <= to_signed(-998,32);
				when 2007 => sin_data_int <= to_signed(63,32); cos_data_int <= to_signed(-998,32);
				when 2008 => sin_data_int <= to_signed(61,32); cos_data_int <= to_signed(-998,32);
				when 2009 => sin_data_int <= to_signed(60,32); cos_data_int <= to_signed(-998,32);
				when 2010 => sin_data_int <= to_signed(58,32); cos_data_int <= to_signed(-998,32);
				when 2011 => sin_data_int <= to_signed(57,32); cos_data_int <= to_signed(-998,32);
				when 2012 => sin_data_int <= to_signed(55,32); cos_data_int <= to_signed(-999,32);
				when 2013 => sin_data_int <= to_signed(54,32); cos_data_int <= to_signed(-999,32);
				when 2014 => sin_data_int <= to_signed(52,32); cos_data_int <= to_signed(-999,32);
				when 2015 => sin_data_int <= to_signed(51,32); cos_data_int <= to_signed(-999,32);
				when 2016 => sin_data_int <= to_signed(49,32); cos_data_int <= to_signed(-999,32);
				when 2017 => sin_data_int <= to_signed(48,32); cos_data_int <= to_signed(-999,32);
				when 2018 => sin_data_int <= to_signed(46,32); cos_data_int <= to_signed(-999,32);
				when 2019 => sin_data_int <= to_signed(44,32); cos_data_int <= to_signed(-999,32);
				when 2020 => sin_data_int <= to_signed(43,32); cos_data_int <= to_signed(-999,32);
				when 2021 => sin_data_int <= to_signed(41,32); cos_data_int <= to_signed(-999,32);
				when 2022 => sin_data_int <= to_signed(40,32); cos_data_int <= to_signed(-999,32);
				when 2023 => sin_data_int <= to_signed(38,32); cos_data_int <= to_signed(-999,32);
				when 2024 => sin_data_int <= to_signed(37,32); cos_data_int <= to_signed(-999,32);
				when 2025 => sin_data_int <= to_signed(35,32); cos_data_int <= to_signed(-999,32);
				when 2026 => sin_data_int <= to_signed(34,32); cos_data_int <= to_signed(-999,32);
				when 2027 => sin_data_int <= to_signed(32,32); cos_data_int <= to_signed(-1000,32);
				when 2028 => sin_data_int <= to_signed(31,32); cos_data_int <= to_signed(-1000,32);
				when 2029 => sin_data_int <= to_signed(29,32); cos_data_int <= to_signed(-1000,32);
				when 2030 => sin_data_int <= to_signed(28,32); cos_data_int <= to_signed(-1000,32);
				when 2031 => sin_data_int <= to_signed(26,32); cos_data_int <= to_signed(-1000,32);
				when 2032 => sin_data_int <= to_signed(25,32); cos_data_int <= to_signed(-1000,32);
				when 2033 => sin_data_int <= to_signed(23,32); cos_data_int <= to_signed(-1000,32);
				when 2034 => sin_data_int <= to_signed(21,32); cos_data_int <= to_signed(-1000,32);
				when 2035 => sin_data_int <= to_signed(20,32); cos_data_int <= to_signed(-1000,32);
				when 2036 => sin_data_int <= to_signed(18,32); cos_data_int <= to_signed(-1000,32);
				when 2037 => sin_data_int <= to_signed(17,32); cos_data_int <= to_signed(-1000,32);
				when 2038 => sin_data_int <= to_signed(15,32); cos_data_int <= to_signed(-1000,32);
				when 2039 => sin_data_int <= to_signed(14,32); cos_data_int <= to_signed(-1000,32);
				when 2040 => sin_data_int <= to_signed(12,32); cos_data_int <= to_signed(-1000,32);
				when 2041 => sin_data_int <= to_signed(11,32); cos_data_int <= to_signed(-1000,32);
				when 2042 => sin_data_int <= to_signed(9,32); cos_data_int <= to_signed(-1000,32);
				when 2043 => sin_data_int <= to_signed(8,32); cos_data_int <= to_signed(-1000,32);
				when 2044 => sin_data_int <= to_signed(6,32); cos_data_int <= to_signed(-1000,32);
				when 2045 => sin_data_int <= to_signed(5,32); cos_data_int <= to_signed(-1000,32);
				when 2046 => sin_data_int <= to_signed(3,32); cos_data_int <= to_signed(-1000,32);
				when 2047 => sin_data_int <= to_signed(2,32); cos_data_int <= to_signed(-1000,32);
				when 2048 => sin_data_int <= to_signed(0,32); cos_data_int <= to_signed(-1000,32);
				when 2049 => sin_data_int <= to_signed(-2,32); cos_data_int <= to_signed(-1000,32);
				when 2050 => sin_data_int <= to_signed(-3,32); cos_data_int <= to_signed(-1000,32);
				when 2051 => sin_data_int <= to_signed(-5,32); cos_data_int <= to_signed(-1000,32);
				when 2052 => sin_data_int <= to_signed(-6,32); cos_data_int <= to_signed(-1000,32);
				when 2053 => sin_data_int <= to_signed(-8,32); cos_data_int <= to_signed(-1000,32);
				when 2054 => sin_data_int <= to_signed(-9,32); cos_data_int <= to_signed(-1000,32);
				when 2055 => sin_data_int <= to_signed(-11,32); cos_data_int <= to_signed(-1000,32);
				when 2056 => sin_data_int <= to_signed(-12,32); cos_data_int <= to_signed(-1000,32);
				when 2057 => sin_data_int <= to_signed(-14,32); cos_data_int <= to_signed(-1000,32);
				when 2058 => sin_data_int <= to_signed(-15,32); cos_data_int <= to_signed(-1000,32);
				when 2059 => sin_data_int <= to_signed(-17,32); cos_data_int <= to_signed(-1000,32);
				when 2060 => sin_data_int <= to_signed(-18,32); cos_data_int <= to_signed(-1000,32);
				when 2061 => sin_data_int <= to_signed(-20,32); cos_data_int <= to_signed(-1000,32);
				when 2062 => sin_data_int <= to_signed(-21,32); cos_data_int <= to_signed(-1000,32);
				when 2063 => sin_data_int <= to_signed(-23,32); cos_data_int <= to_signed(-1000,32);
				when 2064 => sin_data_int <= to_signed(-25,32); cos_data_int <= to_signed(-1000,32);
				when 2065 => sin_data_int <= to_signed(-26,32); cos_data_int <= to_signed(-1000,32);
				when 2066 => sin_data_int <= to_signed(-28,32); cos_data_int <= to_signed(-1000,32);
				when 2067 => sin_data_int <= to_signed(-29,32); cos_data_int <= to_signed(-1000,32);
				when 2068 => sin_data_int <= to_signed(-31,32); cos_data_int <= to_signed(-999,32);
				when 2069 => sin_data_int <= to_signed(-32,32); cos_data_int <= to_signed(-999,32);
				when 2070 => sin_data_int <= to_signed(-34,32); cos_data_int <= to_signed(-999,32);
				when 2071 => sin_data_int <= to_signed(-35,32); cos_data_int <= to_signed(-999,32);
				when 2072 => sin_data_int <= to_signed(-37,32); cos_data_int <= to_signed(-999,32);
				when 2073 => sin_data_int <= to_signed(-38,32); cos_data_int <= to_signed(-999,32);
				when 2074 => sin_data_int <= to_signed(-40,32); cos_data_int <= to_signed(-999,32);
				when 2075 => sin_data_int <= to_signed(-41,32); cos_data_int <= to_signed(-999,32);
				when 2076 => sin_data_int <= to_signed(-43,32); cos_data_int <= to_signed(-999,32);
				when 2077 => sin_data_int <= to_signed(-44,32); cos_data_int <= to_signed(-999,32);
				when 2078 => sin_data_int <= to_signed(-46,32); cos_data_int <= to_signed(-999,32);
				when 2079 => sin_data_int <= to_signed(-48,32); cos_data_int <= to_signed(-999,32);
				when 2080 => sin_data_int <= to_signed(-49,32); cos_data_int <= to_signed(-999,32);
				when 2081 => sin_data_int <= to_signed(-51,32); cos_data_int <= to_signed(-999,32);
				when 2082 => sin_data_int <= to_signed(-52,32); cos_data_int <= to_signed(-999,32);
				when 2083 => sin_data_int <= to_signed(-54,32); cos_data_int <= to_signed(-998,32);
				when 2084 => sin_data_int <= to_signed(-55,32); cos_data_int <= to_signed(-998,32);
				when 2085 => sin_data_int <= to_signed(-57,32); cos_data_int <= to_signed(-998,32);
				when 2086 => sin_data_int <= to_signed(-58,32); cos_data_int <= to_signed(-998,32);
				when 2087 => sin_data_int <= to_signed(-60,32); cos_data_int <= to_signed(-998,32);
				when 2088 => sin_data_int <= to_signed(-61,32); cos_data_int <= to_signed(-998,32);
				when 2089 => sin_data_int <= to_signed(-63,32); cos_data_int <= to_signed(-998,32);
				when 2090 => sin_data_int <= to_signed(-64,32); cos_data_int <= to_signed(-998,32);
				when 2091 => sin_data_int <= to_signed(-66,32); cos_data_int <= to_signed(-998,32);
				when 2092 => sin_data_int <= to_signed(-67,32); cos_data_int <= to_signed(-998,32);
				when 2093 => sin_data_int <= to_signed(-69,32); cos_data_int <= to_signed(-998,32);
				when 2094 => sin_data_int <= to_signed(-71,32); cos_data_int <= to_signed(-997,32);
				when 2095 => sin_data_int <= to_signed(-72,32); cos_data_int <= to_signed(-997,32);
				when 2096 => sin_data_int <= to_signed(-74,32); cos_data_int <= to_signed(-997,32);
				when 2097 => sin_data_int <= to_signed(-75,32); cos_data_int <= to_signed(-997,32);
				when 2098 => sin_data_int <= to_signed(-77,32); cos_data_int <= to_signed(-997,32);
				when 2099 => sin_data_int <= to_signed(-78,32); cos_data_int <= to_signed(-997,32);
				when 2100 => sin_data_int <= to_signed(-80,32); cos_data_int <= to_signed(-997,32);
				when 2101 => sin_data_int <= to_signed(-81,32); cos_data_int <= to_signed(-997,32);
				when 2102 => sin_data_int <= to_signed(-83,32); cos_data_int <= to_signed(-996,32);
				when 2103 => sin_data_int <= to_signed(-84,32); cos_data_int <= to_signed(-996,32);
				when 2104 => sin_data_int <= to_signed(-86,32); cos_data_int <= to_signed(-996,32);
				when 2105 => sin_data_int <= to_signed(-87,32); cos_data_int <= to_signed(-996,32);
				when 2106 => sin_data_int <= to_signed(-89,32); cos_data_int <= to_signed(-996,32);
				when 2107 => sin_data_int <= to_signed(-90,32); cos_data_int <= to_signed(-996,32);
				when 2108 => sin_data_int <= to_signed(-92,32); cos_data_int <= to_signed(-996,32);
				when 2109 => sin_data_int <= to_signed(-93,32); cos_data_int <= to_signed(-995,32);
				when 2110 => sin_data_int <= to_signed(-95,32); cos_data_int <= to_signed(-995,32);
				when 2111 => sin_data_int <= to_signed(-96,32); cos_data_int <= to_signed(-995,32);
				when 2112 => sin_data_int <= to_signed(-98,32); cos_data_int <= to_signed(-995,32);
				when 2113 => sin_data_int <= to_signed(-100,32); cos_data_int <= to_signed(-995,32);
				when 2114 => sin_data_int <= to_signed(-101,32); cos_data_int <= to_signed(-995,32);
				when 2115 => sin_data_int <= to_signed(-103,32); cos_data_int <= to_signed(-995,32);
				when 2116 => sin_data_int <= to_signed(-104,32); cos_data_int <= to_signed(-994,32);
				when 2117 => sin_data_int <= to_signed(-106,32); cos_data_int <= to_signed(-994,32);
				when 2118 => sin_data_int <= to_signed(-107,32); cos_data_int <= to_signed(-994,32);
				when 2119 => sin_data_int <= to_signed(-109,32); cos_data_int <= to_signed(-994,32);
				when 2120 => sin_data_int <= to_signed(-110,32); cos_data_int <= to_signed(-994,32);
				when 2121 => sin_data_int <= to_signed(-112,32); cos_data_int <= to_signed(-994,32);
				when 2122 => sin_data_int <= to_signed(-113,32); cos_data_int <= to_signed(-993,32);
				when 2123 => sin_data_int <= to_signed(-115,32); cos_data_int <= to_signed(-993,32);
				when 2124 => sin_data_int <= to_signed(-116,32); cos_data_int <= to_signed(-993,32);
				when 2125 => sin_data_int <= to_signed(-118,32); cos_data_int <= to_signed(-993,32);
				when 2126 => sin_data_int <= to_signed(-119,32); cos_data_int <= to_signed(-993,32);
				when 2127 => sin_data_int <= to_signed(-121,32); cos_data_int <= to_signed(-992,32);
				when 2128 => sin_data_int <= to_signed(-122,32); cos_data_int <= to_signed(-992,32);
				when 2129 => sin_data_int <= to_signed(-124,32); cos_data_int <= to_signed(-992,32);
				when 2130 => sin_data_int <= to_signed(-125,32); cos_data_int <= to_signed(-992,32);
				when 2131 => sin_data_int <= to_signed(-127,32); cos_data_int <= to_signed(-992,32);
				when 2132 => sin_data_int <= to_signed(-128,32); cos_data_int <= to_signed(-992,32);
				when 2133 => sin_data_int <= to_signed(-130,32); cos_data_int <= to_signed(-991,32);
				when 2134 => sin_data_int <= to_signed(-132,32); cos_data_int <= to_signed(-991,32);
				when 2135 => sin_data_int <= to_signed(-133,32); cos_data_int <= to_signed(-991,32);
				when 2136 => sin_data_int <= to_signed(-135,32); cos_data_int <= to_signed(-991,32);
				when 2137 => sin_data_int <= to_signed(-136,32); cos_data_int <= to_signed(-990,32);
				when 2138 => sin_data_int <= to_signed(-138,32); cos_data_int <= to_signed(-990,32);
				when 2139 => sin_data_int <= to_signed(-139,32); cos_data_int <= to_signed(-990,32);
				when 2140 => sin_data_int <= to_signed(-141,32); cos_data_int <= to_signed(-990,32);
				when 2141 => sin_data_int <= to_signed(-142,32); cos_data_int <= to_signed(-990,32);
				when 2142 => sin_data_int <= to_signed(-144,32); cos_data_int <= to_signed(-989,32);
				when 2143 => sin_data_int <= to_signed(-145,32); cos_data_int <= to_signed(-989,32);
				when 2144 => sin_data_int <= to_signed(-147,32); cos_data_int <= to_signed(-989,32);
				when 2145 => sin_data_int <= to_signed(-148,32); cos_data_int <= to_signed(-989,32);
				when 2146 => sin_data_int <= to_signed(-150,32); cos_data_int <= to_signed(-988,32);
				when 2147 => sin_data_int <= to_signed(-151,32); cos_data_int <= to_signed(-988,32);
				when 2148 => sin_data_int <= to_signed(-153,32); cos_data_int <= to_signed(-988,32);
				when 2149 => sin_data_int <= to_signed(-154,32); cos_data_int <= to_signed(-988,32);
				when 2150 => sin_data_int <= to_signed(-156,32); cos_data_int <= to_signed(-988,32);
				when 2151 => sin_data_int <= to_signed(-157,32); cos_data_int <= to_signed(-987,32);
				when 2152 => sin_data_int <= to_signed(-159,32); cos_data_int <= to_signed(-987,32);
				when 2153 => sin_data_int <= to_signed(-160,32); cos_data_int <= to_signed(-987,32);
				when 2154 => sin_data_int <= to_signed(-162,32); cos_data_int <= to_signed(-987,32);
				when 2155 => sin_data_int <= to_signed(-163,32); cos_data_int <= to_signed(-986,32);
				when 2156 => sin_data_int <= to_signed(-165,32); cos_data_int <= to_signed(-986,32);
				when 2157 => sin_data_int <= to_signed(-166,32); cos_data_int <= to_signed(-986,32);
				when 2158 => sin_data_int <= to_signed(-168,32); cos_data_int <= to_signed(-986,32);
				when 2159 => sin_data_int <= to_signed(-169,32); cos_data_int <= to_signed(-985,32);
				when 2160 => sin_data_int <= to_signed(-171,32); cos_data_int <= to_signed(-985,32);
				when 2161 => sin_data_int <= to_signed(-172,32); cos_data_int <= to_signed(-985,32);
				when 2162 => sin_data_int <= to_signed(-174,32); cos_data_int <= to_signed(-984,32);
				when 2163 => sin_data_int <= to_signed(-175,32); cos_data_int <= to_signed(-984,32);
				when 2164 => sin_data_int <= to_signed(-177,32); cos_data_int <= to_signed(-984,32);
				when 2165 => sin_data_int <= to_signed(-179,32); cos_data_int <= to_signed(-984,32);
				when 2166 => sin_data_int <= to_signed(-180,32); cos_data_int <= to_signed(-983,32);
				when 2167 => sin_data_int <= to_signed(-182,32); cos_data_int <= to_signed(-983,32);
				when 2168 => sin_data_int <= to_signed(-183,32); cos_data_int <= to_signed(-983,32);
				when 2169 => sin_data_int <= to_signed(-185,32); cos_data_int <= to_signed(-983,32);
				when 2170 => sin_data_int <= to_signed(-186,32); cos_data_int <= to_signed(-982,32);
				when 2171 => sin_data_int <= to_signed(-188,32); cos_data_int <= to_signed(-982,32);
				when 2172 => sin_data_int <= to_signed(-189,32); cos_data_int <= to_signed(-982,32);
				when 2173 => sin_data_int <= to_signed(-191,32); cos_data_int <= to_signed(-981,32);
				when 2174 => sin_data_int <= to_signed(-192,32); cos_data_int <= to_signed(-981,32);
				when 2175 => sin_data_int <= to_signed(-194,32); cos_data_int <= to_signed(-981,32);
				when 2176 => sin_data_int <= to_signed(-195,32); cos_data_int <= to_signed(-980,32);
				when 2177 => sin_data_int <= to_signed(-197,32); cos_data_int <= to_signed(-980,32);
				when 2178 => sin_data_int <= to_signed(-198,32); cos_data_int <= to_signed(-980,32);
				when 2179 => sin_data_int <= to_signed(-200,32); cos_data_int <= to_signed(-980,32);
				when 2180 => sin_data_int <= to_signed(-201,32); cos_data_int <= to_signed(-979,32);
				when 2181 => sin_data_int <= to_signed(-203,32); cos_data_int <= to_signed(-979,32);
				when 2182 => sin_data_int <= to_signed(-204,32); cos_data_int <= to_signed(-979,32);
				when 2183 => sin_data_int <= to_signed(-206,32); cos_data_int <= to_signed(-978,32);
				when 2184 => sin_data_int <= to_signed(-207,32); cos_data_int <= to_signed(-978,32);
				when 2185 => sin_data_int <= to_signed(-209,32); cos_data_int <= to_signed(-978,32);
				when 2186 => sin_data_int <= to_signed(-210,32); cos_data_int <= to_signed(-977,32);
				when 2187 => sin_data_int <= to_signed(-212,32); cos_data_int <= to_signed(-977,32);
				when 2188 => sin_data_int <= to_signed(-213,32); cos_data_int <= to_signed(-977,32);
				when 2189 => sin_data_int <= to_signed(-215,32); cos_data_int <= to_signed(-976,32);
				when 2190 => sin_data_int <= to_signed(-216,32); cos_data_int <= to_signed(-976,32);
				when 2191 => sin_data_int <= to_signed(-218,32); cos_data_int <= to_signed(-976,32);
				when 2192 => sin_data_int <= to_signed(-219,32); cos_data_int <= to_signed(-975,32);
				when 2193 => sin_data_int <= to_signed(-221,32); cos_data_int <= to_signed(-975,32);
				when 2194 => sin_data_int <= to_signed(-222,32); cos_data_int <= to_signed(-975,32);
				when 2195 => sin_data_int <= to_signed(-224,32); cos_data_int <= to_signed(-974,32);
				when 2196 => sin_data_int <= to_signed(-225,32); cos_data_int <= to_signed(-974,32);
				when 2197 => sin_data_int <= to_signed(-227,32); cos_data_int <= to_signed(-974,32);
				when 2198 => sin_data_int <= to_signed(-228,32); cos_data_int <= to_signed(-973,32);
				when 2199 => sin_data_int <= to_signed(-230,32); cos_data_int <= to_signed(-973,32);
				when 2200 => sin_data_int <= to_signed(-231,32); cos_data_int <= to_signed(-973,32);
				when 2201 => sin_data_int <= to_signed(-233,32); cos_data_int <= to_signed(-972,32);
				when 2202 => sin_data_int <= to_signed(-234,32); cos_data_int <= to_signed(-972,32);
				when 2203 => sin_data_int <= to_signed(-236,32); cos_data_int <= to_signed(-972,32);
				when 2204 => sin_data_int <= to_signed(-237,32); cos_data_int <= to_signed(-971,32);
				when 2205 => sin_data_int <= to_signed(-239,32); cos_data_int <= to_signed(-971,32);
				when 2206 => sin_data_int <= to_signed(-240,32); cos_data_int <= to_signed(-970,32);
				when 2207 => sin_data_int <= to_signed(-241,32); cos_data_int <= to_signed(-970,32);
				when 2208 => sin_data_int <= to_signed(-243,32); cos_data_int <= to_signed(-970,32);
				when 2209 => sin_data_int <= to_signed(-244,32); cos_data_int <= to_signed(-969,32);
				when 2210 => sin_data_int <= to_signed(-246,32); cos_data_int <= to_signed(-969,32);
				when 2211 => sin_data_int <= to_signed(-247,32); cos_data_int <= to_signed(-969,32);
				when 2212 => sin_data_int <= to_signed(-249,32); cos_data_int <= to_signed(-968,32);
				when 2213 => sin_data_int <= to_signed(-250,32); cos_data_int <= to_signed(-968,32);
				when 2214 => sin_data_int <= to_signed(-252,32); cos_data_int <= to_signed(-967,32);
				when 2215 => sin_data_int <= to_signed(-253,32); cos_data_int <= to_signed(-967,32);
				when 2216 => sin_data_int <= to_signed(-255,32); cos_data_int <= to_signed(-967,32);
				when 2217 => sin_data_int <= to_signed(-256,32); cos_data_int <= to_signed(-966,32);
				when 2218 => sin_data_int <= to_signed(-258,32); cos_data_int <= to_signed(-966,32);
				when 2219 => sin_data_int <= to_signed(-259,32); cos_data_int <= to_signed(-965,32);
				when 2220 => sin_data_int <= to_signed(-261,32); cos_data_int <= to_signed(-965,32);
				when 2221 => sin_data_int <= to_signed(-262,32); cos_data_int <= to_signed(-965,32);
				when 2222 => sin_data_int <= to_signed(-264,32); cos_data_int <= to_signed(-964,32);
				when 2223 => sin_data_int <= to_signed(-265,32); cos_data_int <= to_signed(-964,32);
				when 2224 => sin_data_int <= to_signed(-267,32); cos_data_int <= to_signed(-963,32);
				when 2225 => sin_data_int <= to_signed(-268,32); cos_data_int <= to_signed(-963,32);
				when 2226 => sin_data_int <= to_signed(-270,32); cos_data_int <= to_signed(-963,32);
				when 2227 => sin_data_int <= to_signed(-271,32); cos_data_int <= to_signed(-962,32);
				when 2228 => sin_data_int <= to_signed(-273,32); cos_data_int <= to_signed(-962,32);
				when 2229 => sin_data_int <= to_signed(-274,32); cos_data_int <= to_signed(-961,32);
				when 2230 => sin_data_int <= to_signed(-276,32); cos_data_int <= to_signed(-961,32);
				when 2231 => sin_data_int <= to_signed(-277,32); cos_data_int <= to_signed(-960,32);
				when 2232 => sin_data_int <= to_signed(-279,32); cos_data_int <= to_signed(-960,32);
				when 2233 => sin_data_int <= to_signed(-280,32); cos_data_int <= to_signed(-960,32);
				when 2234 => sin_data_int <= to_signed(-281,32); cos_data_int <= to_signed(-959,32);
				when 2235 => sin_data_int <= to_signed(-283,32); cos_data_int <= to_signed(-959,32);
				when 2236 => sin_data_int <= to_signed(-284,32); cos_data_int <= to_signed(-958,32);
				when 2237 => sin_data_int <= to_signed(-286,32); cos_data_int <= to_signed(-958,32);
				when 2238 => sin_data_int <= to_signed(-287,32); cos_data_int <= to_signed(-957,32);
				when 2239 => sin_data_int <= to_signed(-289,32); cos_data_int <= to_signed(-957,32);
				when 2240 => sin_data_int <= to_signed(-290,32); cos_data_int <= to_signed(-956,32);
				when 2241 => sin_data_int <= to_signed(-292,32); cos_data_int <= to_signed(-956,32);
				when 2242 => sin_data_int <= to_signed(-293,32); cos_data_int <= to_signed(-956,32);
				when 2243 => sin_data_int <= to_signed(-295,32); cos_data_int <= to_signed(-955,32);
				when 2244 => sin_data_int <= to_signed(-296,32); cos_data_int <= to_signed(-955,32);
				when 2245 => sin_data_int <= to_signed(-298,32); cos_data_int <= to_signed(-954,32);
				when 2246 => sin_data_int <= to_signed(-299,32); cos_data_int <= to_signed(-954,32);
				when 2247 => sin_data_int <= to_signed(-301,32); cos_data_int <= to_signed(-953,32);
				when 2248 => sin_data_int <= to_signed(-302,32); cos_data_int <= to_signed(-953,32);
				when 2249 => sin_data_int <= to_signed(-303,32); cos_data_int <= to_signed(-952,32);
				when 2250 => sin_data_int <= to_signed(-305,32); cos_data_int <= to_signed(-952,32);
				when 2251 => sin_data_int <= to_signed(-306,32); cos_data_int <= to_signed(-951,32);
				when 2252 => sin_data_int <= to_signed(-308,32); cos_data_int <= to_signed(-951,32);
				when 2253 => sin_data_int <= to_signed(-309,32); cos_data_int <= to_signed(-950,32);
				when 2254 => sin_data_int <= to_signed(-311,32); cos_data_int <= to_signed(-950,32);
				when 2255 => sin_data_int <= to_signed(-312,32); cos_data_int <= to_signed(-950,32);
				when 2256 => sin_data_int <= to_signed(-314,32); cos_data_int <= to_signed(-949,32);
				when 2257 => sin_data_int <= to_signed(-315,32); cos_data_int <= to_signed(-949,32);
				when 2258 => sin_data_int <= to_signed(-317,32); cos_data_int <= to_signed(-948,32);
				when 2259 => sin_data_int <= to_signed(-318,32); cos_data_int <= to_signed(-948,32);
				when 2260 => sin_data_int <= to_signed(-320,32); cos_data_int <= to_signed(-947,32);
				when 2261 => sin_data_int <= to_signed(-321,32); cos_data_int <= to_signed(-947,32);
				when 2262 => sin_data_int <= to_signed(-322,32); cos_data_int <= to_signed(-946,32);
				when 2263 => sin_data_int <= to_signed(-324,32); cos_data_int <= to_signed(-946,32);
				when 2264 => sin_data_int <= to_signed(-325,32); cos_data_int <= to_signed(-945,32);
				when 2265 => sin_data_int <= to_signed(-327,32); cos_data_int <= to_signed(-945,32);
				when 2266 => sin_data_int <= to_signed(-328,32); cos_data_int <= to_signed(-944,32);
				when 2267 => sin_data_int <= to_signed(-330,32); cos_data_int <= to_signed(-944,32);
				when 2268 => sin_data_int <= to_signed(-331,32); cos_data_int <= to_signed(-943,32);
				when 2269 => sin_data_int <= to_signed(-333,32); cos_data_int <= to_signed(-943,32);
				when 2270 => sin_data_int <= to_signed(-334,32); cos_data_int <= to_signed(-942,32);
				when 2271 => sin_data_int <= to_signed(-335,32); cos_data_int <= to_signed(-942,32);
				when 2272 => sin_data_int <= to_signed(-337,32); cos_data_int <= to_signed(-941,32);
				when 2273 => sin_data_int <= to_signed(-338,32); cos_data_int <= to_signed(-941,32);
				when 2274 => sin_data_int <= to_signed(-340,32); cos_data_int <= to_signed(-940,32);
				when 2275 => sin_data_int <= to_signed(-341,32); cos_data_int <= to_signed(-939,32);
				when 2276 => sin_data_int <= to_signed(-343,32); cos_data_int <= to_signed(-939,32);
				when 2277 => sin_data_int <= to_signed(-344,32); cos_data_int <= to_signed(-938,32);
				when 2278 => sin_data_int <= to_signed(-346,32); cos_data_int <= to_signed(-938,32);
				when 2279 => sin_data_int <= to_signed(-347,32); cos_data_int <= to_signed(-937,32);
				when 2280 => sin_data_int <= to_signed(-348,32); cos_data_int <= to_signed(-937,32);
				when 2281 => sin_data_int <= to_signed(-350,32); cos_data_int <= to_signed(-936,32);
				when 2282 => sin_data_int <= to_signed(-351,32); cos_data_int <= to_signed(-936,32);
				when 2283 => sin_data_int <= to_signed(-353,32); cos_data_int <= to_signed(-935,32);
				when 2284 => sin_data_int <= to_signed(-354,32); cos_data_int <= to_signed(-935,32);
				when 2285 => sin_data_int <= to_signed(-356,32); cos_data_int <= to_signed(-934,32);
				when 2286 => sin_data_int <= to_signed(-357,32); cos_data_int <= to_signed(-934,32);
				when 2287 => sin_data_int <= to_signed(-358,32); cos_data_int <= to_signed(-933,32);
				when 2288 => sin_data_int <= to_signed(-360,32); cos_data_int <= to_signed(-932,32);
				when 2289 => sin_data_int <= to_signed(-361,32); cos_data_int <= to_signed(-932,32);
				when 2290 => sin_data_int <= to_signed(-363,32); cos_data_int <= to_signed(-931,32);
				when 2291 => sin_data_int <= to_signed(-364,32); cos_data_int <= to_signed(-931,32);
				when 2292 => sin_data_int <= to_signed(-366,32); cos_data_int <= to_signed(-930,32);
				when 2293 => sin_data_int <= to_signed(-367,32); cos_data_int <= to_signed(-930,32);
				when 2294 => sin_data_int <= to_signed(-368,32); cos_data_int <= to_signed(-929,32);
				when 2295 => sin_data_int <= to_signed(-370,32); cos_data_int <= to_signed(-929,32);
				when 2296 => sin_data_int <= to_signed(-371,32); cos_data_int <= to_signed(-928,32);
				when 2297 => sin_data_int <= to_signed(-373,32); cos_data_int <= to_signed(-927,32);
				when 2298 => sin_data_int <= to_signed(-374,32); cos_data_int <= to_signed(-927,32);
				when 2299 => sin_data_int <= to_signed(-376,32); cos_data_int <= to_signed(-926,32);
				when 2300 => sin_data_int <= to_signed(-377,32); cos_data_int <= to_signed(-926,32);
				when 2301 => sin_data_int <= to_signed(-378,32); cos_data_int <= to_signed(-925,32);
				when 2302 => sin_data_int <= to_signed(-380,32); cos_data_int <= to_signed(-924,32);
				when 2303 => sin_data_int <= to_signed(-381,32); cos_data_int <= to_signed(-924,32);
				when 2304 => sin_data_int <= to_signed(-383,32); cos_data_int <= to_signed(-923,32);
				when 2305 => sin_data_int <= to_signed(-384,32); cos_data_int <= to_signed(-923,32);
				when 2306 => sin_data_int <= to_signed(-386,32); cos_data_int <= to_signed(-922,32);
				when 2307 => sin_data_int <= to_signed(-387,32); cos_data_int <= to_signed(-922,32);
				when 2308 => sin_data_int <= to_signed(-388,32); cos_data_int <= to_signed(-921,32);
				when 2309 => sin_data_int <= to_signed(-390,32); cos_data_int <= to_signed(-920,32);
				when 2310 => sin_data_int <= to_signed(-391,32); cos_data_int <= to_signed(-920,32);
				when 2311 => sin_data_int <= to_signed(-393,32); cos_data_int <= to_signed(-919,32);
				when 2312 => sin_data_int <= to_signed(-394,32); cos_data_int <= to_signed(-919,32);
				when 2313 => sin_data_int <= to_signed(-395,32); cos_data_int <= to_signed(-918,32);
				when 2314 => sin_data_int <= to_signed(-397,32); cos_data_int <= to_signed(-917,32);
				when 2315 => sin_data_int <= to_signed(-398,32); cos_data_int <= to_signed(-917,32);
				when 2316 => sin_data_int <= to_signed(-400,32); cos_data_int <= to_signed(-916,32);
				when 2317 => sin_data_int <= to_signed(-401,32); cos_data_int <= to_signed(-915,32);
				when 2318 => sin_data_int <= to_signed(-402,32); cos_data_int <= to_signed(-915,32);
				when 2319 => sin_data_int <= to_signed(-404,32); cos_data_int <= to_signed(-914,32);
				when 2320 => sin_data_int <= to_signed(-405,32); cos_data_int <= to_signed(-914,32);
				when 2321 => sin_data_int <= to_signed(-407,32); cos_data_int <= to_signed(-913,32);
				when 2322 => sin_data_int <= to_signed(-408,32); cos_data_int <= to_signed(-912,32);
				when 2323 => sin_data_int <= to_signed(-409,32); cos_data_int <= to_signed(-912,32);
				when 2324 => sin_data_int <= to_signed(-411,32); cos_data_int <= to_signed(-911,32);
				when 2325 => sin_data_int <= to_signed(-412,32); cos_data_int <= to_signed(-910,32);
				when 2326 => sin_data_int <= to_signed(-414,32); cos_data_int <= to_signed(-910,32);
				when 2327 => sin_data_int <= to_signed(-415,32); cos_data_int <= to_signed(-909,32);
				when 2328 => sin_data_int <= to_signed(-416,32); cos_data_int <= to_signed(-909,32);
				when 2329 => sin_data_int <= to_signed(-418,32); cos_data_int <= to_signed(-908,32);
				when 2330 => sin_data_int <= to_signed(-419,32); cos_data_int <= to_signed(-907,32);
				when 2331 => sin_data_int <= to_signed(-421,32); cos_data_int <= to_signed(-907,32);
				when 2332 => sin_data_int <= to_signed(-422,32); cos_data_int <= to_signed(-906,32);
				when 2333 => sin_data_int <= to_signed(-423,32); cos_data_int <= to_signed(-905,32);
				when 2334 => sin_data_int <= to_signed(-425,32); cos_data_int <= to_signed(-905,32);
				when 2335 => sin_data_int <= to_signed(-426,32); cos_data_int <= to_signed(-904,32);
				when 2336 => sin_data_int <= to_signed(-428,32); cos_data_int <= to_signed(-903,32);
				when 2337 => sin_data_int <= to_signed(-429,32); cos_data_int <= to_signed(-903,32);
				when 2338 => sin_data_int <= to_signed(-430,32); cos_data_int <= to_signed(-902,32);
				when 2339 => sin_data_int <= to_signed(-432,32); cos_data_int <= to_signed(-901,32);
				when 2340 => sin_data_int <= to_signed(-433,32); cos_data_int <= to_signed(-901,32);
				when 2341 => sin_data_int <= to_signed(-434,32); cos_data_int <= to_signed(-900,32);
				when 2342 => sin_data_int <= to_signed(-436,32); cos_data_int <= to_signed(-899,32);
				when 2343 => sin_data_int <= to_signed(-437,32); cos_data_int <= to_signed(-899,32);
				when 2344 => sin_data_int <= to_signed(-439,32); cos_data_int <= to_signed(-898,32);
				when 2345 => sin_data_int <= to_signed(-440,32); cos_data_int <= to_signed(-897,32);
				when 2346 => sin_data_int <= to_signed(-441,32); cos_data_int <= to_signed(-897,32);
				when 2347 => sin_data_int <= to_signed(-443,32); cos_data_int <= to_signed(-896,32);
				when 2348 => sin_data_int <= to_signed(-444,32); cos_data_int <= to_signed(-895,32);
				when 2349 => sin_data_int <= to_signed(-445,32); cos_data_int <= to_signed(-895,32);
				when 2350 => sin_data_int <= to_signed(-447,32); cos_data_int <= to_signed(-894,32);
				when 2351 => sin_data_int <= to_signed(-448,32); cos_data_int <= to_signed(-893,32);
				when 2352 => sin_data_int <= to_signed(-450,32); cos_data_int <= to_signed(-893,32);
				when 2353 => sin_data_int <= to_signed(-451,32); cos_data_int <= to_signed(-892,32);
				when 2354 => sin_data_int <= to_signed(-452,32); cos_data_int <= to_signed(-891,32);
				when 2355 => sin_data_int <= to_signed(-454,32); cos_data_int <= to_signed(-890,32);
				when 2356 => sin_data_int <= to_signed(-455,32); cos_data_int <= to_signed(-890,32);
				when 2357 => sin_data_int <= to_signed(-456,32); cos_data_int <= to_signed(-889,32);
				when 2358 => sin_data_int <= to_signed(-458,32); cos_data_int <= to_signed(-888,32);
				when 2359 => sin_data_int <= to_signed(-459,32); cos_data_int <= to_signed(-888,32);
				when 2360 => sin_data_int <= to_signed(-461,32); cos_data_int <= to_signed(-887,32);
				when 2361 => sin_data_int <= to_signed(-462,32); cos_data_int <= to_signed(-886,32);
				when 2362 => sin_data_int <= to_signed(-463,32); cos_data_int <= to_signed(-886,32);
				when 2363 => sin_data_int <= to_signed(-465,32); cos_data_int <= to_signed(-885,32);
				when 2364 => sin_data_int <= to_signed(-466,32); cos_data_int <= to_signed(-884,32);
				when 2365 => sin_data_int <= to_signed(-467,32); cos_data_int <= to_signed(-883,32);
				when 2366 => sin_data_int <= to_signed(-469,32); cos_data_int <= to_signed(-883,32);
				when 2367 => sin_data_int <= to_signed(-470,32); cos_data_int <= to_signed(-882,32);
				when 2368 => sin_data_int <= to_signed(-471,32); cos_data_int <= to_signed(-881,32);
				when 2369 => sin_data_int <= to_signed(-473,32); cos_data_int <= to_signed(-880,32);
				when 2370 => sin_data_int <= to_signed(-474,32); cos_data_int <= to_signed(-880,32);
				when 2371 => sin_data_int <= to_signed(-475,32); cos_data_int <= to_signed(-879,32);
				when 2372 => sin_data_int <= to_signed(-477,32); cos_data_int <= to_signed(-878,32);
				when 2373 => sin_data_int <= to_signed(-478,32); cos_data_int <= to_signed(-878,32);
				when 2374 => sin_data_int <= to_signed(-479,32); cos_data_int <= to_signed(-877,32);
				when 2375 => sin_data_int <= to_signed(-481,32); cos_data_int <= to_signed(-876,32);
				when 2376 => sin_data_int <= to_signed(-482,32); cos_data_int <= to_signed(-875,32);
				when 2377 => sin_data_int <= to_signed(-484,32); cos_data_int <= to_signed(-875,32);
				when 2378 => sin_data_int <= to_signed(-485,32); cos_data_int <= to_signed(-874,32);
				when 2379 => sin_data_int <= to_signed(-486,32); cos_data_int <= to_signed(-873,32);
				when 2380 => sin_data_int <= to_signed(-488,32); cos_data_int <= to_signed(-872,32);
				when 2381 => sin_data_int <= to_signed(-489,32); cos_data_int <= to_signed(-872,32);
				when 2382 => sin_data_int <= to_signed(-490,32); cos_data_int <= to_signed(-871,32);
				when 2383 => sin_data_int <= to_signed(-492,32); cos_data_int <= to_signed(-870,32);
				when 2384 => sin_data_int <= to_signed(-493,32); cos_data_int <= to_signed(-869,32);
				when 2385 => sin_data_int <= to_signed(-494,32); cos_data_int <= to_signed(-869,32);
				when 2386 => sin_data_int <= to_signed(-496,32); cos_data_int <= to_signed(-868,32);
				when 2387 => sin_data_int <= to_signed(-497,32); cos_data_int <= to_signed(-867,32);
				when 2388 => sin_data_int <= to_signed(-498,32); cos_data_int <= to_signed(-866,32);
				when 2389 => sin_data_int <= to_signed(-500,32); cos_data_int <= to_signed(-866,32);
				when 2390 => sin_data_int <= to_signed(-501,32); cos_data_int <= to_signed(-865,32);
				when 2391 => sin_data_int <= to_signed(-502,32); cos_data_int <= to_signed(-864,32);
				when 2392 => sin_data_int <= to_signed(-504,32); cos_data_int <= to_signed(-863,32);
				when 2393 => sin_data_int <= to_signed(-505,32); cos_data_int <= to_signed(-862,32);
				when 2394 => sin_data_int <= to_signed(-506,32); cos_data_int <= to_signed(-862,32);
				when 2395 => sin_data_int <= to_signed(-508,32); cos_data_int <= to_signed(-861,32);
				when 2396 => sin_data_int <= to_signed(-509,32); cos_data_int <= to_signed(-860,32);
				when 2397 => sin_data_int <= to_signed(-510,32); cos_data_int <= to_signed(-859,32);
				when 2398 => sin_data_int <= to_signed(-511,32); cos_data_int <= to_signed(-859,32);
				when 2399 => sin_data_int <= to_signed(-513,32); cos_data_int <= to_signed(-858,32);
				when 2400 => sin_data_int <= to_signed(-514,32); cos_data_int <= to_signed(-857,32);
				when 2401 => sin_data_int <= to_signed(-515,32); cos_data_int <= to_signed(-856,32);
				when 2402 => sin_data_int <= to_signed(-517,32); cos_data_int <= to_signed(-855,32);
				when 2403 => sin_data_int <= to_signed(-518,32); cos_data_int <= to_signed(-855,32);
				when 2404 => sin_data_int <= to_signed(-519,32); cos_data_int <= to_signed(-854,32);
				when 2405 => sin_data_int <= to_signed(-521,32); cos_data_int <= to_signed(-853,32);
				when 2406 => sin_data_int <= to_signed(-522,32); cos_data_int <= to_signed(-852,32);
				when 2407 => sin_data_int <= to_signed(-523,32); cos_data_int <= to_signed(-851,32);
				when 2408 => sin_data_int <= to_signed(-525,32); cos_data_int <= to_signed(-851,32);
				when 2409 => sin_data_int <= to_signed(-526,32); cos_data_int <= to_signed(-850,32);
				when 2410 => sin_data_int <= to_signed(-527,32); cos_data_int <= to_signed(-849,32);
				when 2411 => sin_data_int <= to_signed(-529,32); cos_data_int <= to_signed(-848,32);
				when 2412 => sin_data_int <= to_signed(-530,32); cos_data_int <= to_signed(-847,32);
				when 2413 => sin_data_int <= to_signed(-531,32); cos_data_int <= to_signed(-846,32);
				when 2414 => sin_data_int <= to_signed(-532,32); cos_data_int <= to_signed(-846,32);
				when 2415 => sin_data_int <= to_signed(-534,32); cos_data_int <= to_signed(-845,32);
				when 2416 => sin_data_int <= to_signed(-535,32); cos_data_int <= to_signed(-844,32);
				when 2417 => sin_data_int <= to_signed(-536,32); cos_data_int <= to_signed(-843,32);
				when 2418 => sin_data_int <= to_signed(-538,32); cos_data_int <= to_signed(-842,32);
				when 2419 => sin_data_int <= to_signed(-539,32); cos_data_int <= to_signed(-842,32);
				when 2420 => sin_data_int <= to_signed(-540,32); cos_data_int <= to_signed(-841,32);
				when 2421 => sin_data_int <= to_signed(-541,32); cos_data_int <= to_signed(-840,32);
				when 2422 => sin_data_int <= to_signed(-543,32); cos_data_int <= to_signed(-839,32);
				when 2423 => sin_data_int <= to_signed(-544,32); cos_data_int <= to_signed(-838,32);
				when 2424 => sin_data_int <= to_signed(-545,32); cos_data_int <= to_signed(-837,32);
				when 2425 => sin_data_int <= to_signed(-547,32); cos_data_int <= to_signed(-837,32);
				when 2426 => sin_data_int <= to_signed(-548,32); cos_data_int <= to_signed(-836,32);
				when 2427 => sin_data_int <= to_signed(-549,32); cos_data_int <= to_signed(-835,32);
				when 2428 => sin_data_int <= to_signed(-550,32); cos_data_int <= to_signed(-834,32);
				when 2429 => sin_data_int <= to_signed(-552,32); cos_data_int <= to_signed(-833,32);
				when 2430 => sin_data_int <= to_signed(-553,32); cos_data_int <= to_signed(-832,32);
				when 2431 => sin_data_int <= to_signed(-554,32); cos_data_int <= to_signed(-831,32);
				when 2432 => sin_data_int <= to_signed(-556,32); cos_data_int <= to_signed(-831,32);
				when 2433 => sin_data_int <= to_signed(-557,32); cos_data_int <= to_signed(-830,32);
				when 2434 => sin_data_int <= to_signed(-558,32); cos_data_int <= to_signed(-829,32);
				when 2435 => sin_data_int <= to_signed(-559,32); cos_data_int <= to_signed(-828,32);
				when 2436 => sin_data_int <= to_signed(-561,32); cos_data_int <= to_signed(-827,32);
				when 2437 => sin_data_int <= to_signed(-562,32); cos_data_int <= to_signed(-826,32);
				when 2438 => sin_data_int <= to_signed(-563,32); cos_data_int <= to_signed(-825,32);
				when 2439 => sin_data_int <= to_signed(-564,32); cos_data_int <= to_signed(-825,32);
				when 2440 => sin_data_int <= to_signed(-566,32); cos_data_int <= to_signed(-824,32);
				when 2441 => sin_data_int <= to_signed(-567,32); cos_data_int <= to_signed(-823,32);
				when 2442 => sin_data_int <= to_signed(-568,32); cos_data_int <= to_signed(-822,32);
				when 2443 => sin_data_int <= to_signed(-570,32); cos_data_int <= to_signed(-821,32);
				when 2444 => sin_data_int <= to_signed(-571,32); cos_data_int <= to_signed(-820,32);
				when 2445 => sin_data_int <= to_signed(-572,32); cos_data_int <= to_signed(-819,32);
				when 2446 => sin_data_int <= to_signed(-573,32); cos_data_int <= to_signed(-818,32);
				when 2447 => sin_data_int <= to_signed(-575,32); cos_data_int <= to_signed(-818,32);
				when 2448 => sin_data_int <= to_signed(-576,32); cos_data_int <= to_signed(-817,32);
				when 2449 => sin_data_int <= to_signed(-577,32); cos_data_int <= to_signed(-816,32);
				when 2450 => sin_data_int <= to_signed(-578,32); cos_data_int <= to_signed(-815,32);
				when 2451 => sin_data_int <= to_signed(-580,32); cos_data_int <= to_signed(-814,32);
				when 2452 => sin_data_int <= to_signed(-581,32); cos_data_int <= to_signed(-813,32);
				when 2453 => sin_data_int <= to_signed(-582,32); cos_data_int <= to_signed(-812,32);
				when 2454 => sin_data_int <= to_signed(-583,32); cos_data_int <= to_signed(-811,32);
				when 2455 => sin_data_int <= to_signed(-585,32); cos_data_int <= to_signed(-810,32);
				when 2456 => sin_data_int <= to_signed(-586,32); cos_data_int <= to_signed(-810,32);
				when 2457 => sin_data_int <= to_signed(-587,32); cos_data_int <= to_signed(-809,32);
				when 2458 => sin_data_int <= to_signed(-588,32); cos_data_int <= to_signed(-808,32);
				when 2459 => sin_data_int <= to_signed(-590,32); cos_data_int <= to_signed(-807,32);
				when 2460 => sin_data_int <= to_signed(-591,32); cos_data_int <= to_signed(-806,32);
				when 2461 => sin_data_int <= to_signed(-592,32); cos_data_int <= to_signed(-805,32);
				when 2462 => sin_data_int <= to_signed(-593,32); cos_data_int <= to_signed(-804,32);
				when 2463 => sin_data_int <= to_signed(-594,32); cos_data_int <= to_signed(-803,32);
				when 2464 => sin_data_int <= to_signed(-596,32); cos_data_int <= to_signed(-802,32);
				when 2465 => sin_data_int <= to_signed(-597,32); cos_data_int <= to_signed(-801,32);
				when 2466 => sin_data_int <= to_signed(-598,32); cos_data_int <= to_signed(-800,32);
				when 2467 => sin_data_int <= to_signed(-599,32); cos_data_int <= to_signed(-800,32);
				when 2468 => sin_data_int <= to_signed(-601,32); cos_data_int <= to_signed(-799,32);
				when 2469 => sin_data_int <= to_signed(-602,32); cos_data_int <= to_signed(-798,32);
				when 2470 => sin_data_int <= to_signed(-603,32); cos_data_int <= to_signed(-797,32);
				when 2471 => sin_data_int <= to_signed(-604,32); cos_data_int <= to_signed(-796,32);
				when 2472 => sin_data_int <= to_signed(-606,32); cos_data_int <= to_signed(-795,32);
				when 2473 => sin_data_int <= to_signed(-607,32); cos_data_int <= to_signed(-794,32);
				when 2474 => sin_data_int <= to_signed(-608,32); cos_data_int <= to_signed(-793,32);
				when 2475 => sin_data_int <= to_signed(-609,32); cos_data_int <= to_signed(-792,32);
				when 2476 => sin_data_int <= to_signed(-610,32); cos_data_int <= to_signed(-791,32);
				when 2477 => sin_data_int <= to_signed(-612,32); cos_data_int <= to_signed(-790,32);
				when 2478 => sin_data_int <= to_signed(-613,32); cos_data_int <= to_signed(-789,32);
				when 2479 => sin_data_int <= to_signed(-614,32); cos_data_int <= to_signed(-788,32);
				when 2480 => sin_data_int <= to_signed(-615,32); cos_data_int <= to_signed(-787,32);
				when 2481 => sin_data_int <= to_signed(-616,32); cos_data_int <= to_signed(-786,32);
				when 2482 => sin_data_int <= to_signed(-618,32); cos_data_int <= to_signed(-786,32);
				when 2483 => sin_data_int <= to_signed(-619,32); cos_data_int <= to_signed(-785,32);
				when 2484 => sin_data_int <= to_signed(-620,32); cos_data_int <= to_signed(-784,32);
				when 2485 => sin_data_int <= to_signed(-621,32); cos_data_int <= to_signed(-783,32);
				when 2486 => sin_data_int <= to_signed(-622,32); cos_data_int <= to_signed(-782,32);
				when 2487 => sin_data_int <= to_signed(-624,32); cos_data_int <= to_signed(-781,32);
				when 2488 => sin_data_int <= to_signed(-625,32); cos_data_int <= to_signed(-780,32);
				when 2489 => sin_data_int <= to_signed(-626,32); cos_data_int <= to_signed(-779,32);
				when 2490 => sin_data_int <= to_signed(-627,32); cos_data_int <= to_signed(-778,32);
				when 2491 => sin_data_int <= to_signed(-628,32); cos_data_int <= to_signed(-777,32);
				when 2492 => sin_data_int <= to_signed(-630,32); cos_data_int <= to_signed(-776,32);
				when 2493 => sin_data_int <= to_signed(-631,32); cos_data_int <= to_signed(-775,32);
				when 2494 => sin_data_int <= to_signed(-632,32); cos_data_int <= to_signed(-774,32);
				when 2495 => sin_data_int <= to_signed(-633,32); cos_data_int <= to_signed(-773,32);
				when 2496 => sin_data_int <= to_signed(-634,32); cos_data_int <= to_signed(-772,32);
				when 2497 => sin_data_int <= to_signed(-636,32); cos_data_int <= to_signed(-771,32);
				when 2498 => sin_data_int <= to_signed(-637,32); cos_data_int <= to_signed(-770,32);
				when 2499 => sin_data_int <= to_signed(-638,32); cos_data_int <= to_signed(-769,32);
				when 2500 => sin_data_int <= to_signed(-639,32); cos_data_int <= to_signed(-768,32);
				when 2501 => sin_data_int <= to_signed(-640,32); cos_data_int <= to_signed(-767,32);
				when 2502 => sin_data_int <= to_signed(-641,32); cos_data_int <= to_signed(-766,32);
				when 2503 => sin_data_int <= to_signed(-643,32); cos_data_int <= to_signed(-765,32);
				when 2504 => sin_data_int <= to_signed(-644,32); cos_data_int <= to_signed(-764,32);
				when 2505 => sin_data_int <= to_signed(-645,32); cos_data_int <= to_signed(-763,32);
				when 2506 => sin_data_int <= to_signed(-646,32); cos_data_int <= to_signed(-762,32);
				when 2507 => sin_data_int <= to_signed(-647,32); cos_data_int <= to_signed(-761,32);
				when 2508 => sin_data_int <= to_signed(-649,32); cos_data_int <= to_signed(-760,32);
				when 2509 => sin_data_int <= to_signed(-650,32); cos_data_int <= to_signed(-759,32);
				when 2510 => sin_data_int <= to_signed(-651,32); cos_data_int <= to_signed(-758,32);
				when 2511 => sin_data_int <= to_signed(-652,32); cos_data_int <= to_signed(-757,32);
				when 2512 => sin_data_int <= to_signed(-653,32); cos_data_int <= to_signed(-756,32);
				when 2513 => sin_data_int <= to_signed(-654,32); cos_data_int <= to_signed(-755,32);
				when 2514 => sin_data_int <= to_signed(-655,32); cos_data_int <= to_signed(-754,32);
				when 2515 => sin_data_int <= to_signed(-657,32); cos_data_int <= to_signed(-753,32);
				when 2516 => sin_data_int <= to_signed(-658,32); cos_data_int <= to_signed(-752,32);
				when 2517 => sin_data_int <= to_signed(-659,32); cos_data_int <= to_signed(-751,32);
				when 2518 => sin_data_int <= to_signed(-660,32); cos_data_int <= to_signed(-750,32);
				when 2519 => sin_data_int <= to_signed(-661,32); cos_data_int <= to_signed(-749,32);
				when 2520 => sin_data_int <= to_signed(-662,32); cos_data_int <= to_signed(-748,32);
				when 2521 => sin_data_int <= to_signed(-664,32); cos_data_int <= to_signed(-747,32);
				when 2522 => sin_data_int <= to_signed(-665,32); cos_data_int <= to_signed(-746,32);
				when 2523 => sin_data_int <= to_signed(-666,32); cos_data_int <= to_signed(-745,32);
				when 2524 => sin_data_int <= to_signed(-667,32); cos_data_int <= to_signed(-744,32);
				when 2525 => sin_data_int <= to_signed(-668,32); cos_data_int <= to_signed(-743,32);
				when 2526 => sin_data_int <= to_signed(-669,32); cos_data_int <= to_signed(-742,32);
				when 2527 => sin_data_int <= to_signed(-670,32); cos_data_int <= to_signed(-741,32);
				when 2528 => sin_data_int <= to_signed(-672,32); cos_data_int <= to_signed(-740,32);
				when 2529 => sin_data_int <= to_signed(-673,32); cos_data_int <= to_signed(-739,32);
				when 2530 => sin_data_int <= to_signed(-674,32); cos_data_int <= to_signed(-738,32);
				when 2531 => sin_data_int <= to_signed(-675,32); cos_data_int <= to_signed(-737,32);
				when 2532 => sin_data_int <= to_signed(-676,32); cos_data_int <= to_signed(-736,32);
				when 2533 => sin_data_int <= to_signed(-677,32); cos_data_int <= to_signed(-735,32);
				when 2534 => sin_data_int <= to_signed(-678,32); cos_data_int <= to_signed(-734,32);
				when 2535 => sin_data_int <= to_signed(-679,32); cos_data_int <= to_signed(-733,32);
				when 2536 => sin_data_int <= to_signed(-681,32); cos_data_int <= to_signed(-732,32);
				when 2537 => sin_data_int <= to_signed(-682,32); cos_data_int <= to_signed(-731,32);
				when 2538 => sin_data_int <= to_signed(-683,32); cos_data_int <= to_signed(-730,32);
				when 2539 => sin_data_int <= to_signed(-684,32); cos_data_int <= to_signed(-728,32);
				when 2540 => sin_data_int <= to_signed(-685,32); cos_data_int <= to_signed(-727,32);
				when 2541 => sin_data_int <= to_signed(-686,32); cos_data_int <= to_signed(-726,32);
				when 2542 => sin_data_int <= to_signed(-687,32); cos_data_int <= to_signed(-725,32);
				when 2543 => sin_data_int <= to_signed(-688,32); cos_data_int <= to_signed(-724,32);
				when 2544 => sin_data_int <= to_signed(-690,32); cos_data_int <= to_signed(-723,32);
				when 2545 => sin_data_int <= to_signed(-691,32); cos_data_int <= to_signed(-722,32);
				when 2546 => sin_data_int <= to_signed(-692,32); cos_data_int <= to_signed(-721,32);
				when 2547 => sin_data_int <= to_signed(-693,32); cos_data_int <= to_signed(-720,32);
				when 2548 => sin_data_int <= to_signed(-694,32); cos_data_int <= to_signed(-719,32);
				when 2549 => sin_data_int <= to_signed(-695,32); cos_data_int <= to_signed(-718,32);
				when 2550 => sin_data_int <= to_signed(-696,32); cos_data_int <= to_signed(-717,32);
				when 2551 => sin_data_int <= to_signed(-697,32); cos_data_int <= to_signed(-716,32);
				when 2552 => sin_data_int <= to_signed(-698,32); cos_data_int <= to_signed(-715,32);
				when 2553 => sin_data_int <= to_signed(-699,32); cos_data_int <= to_signed(-714,32);
				when 2554 => sin_data_int <= to_signed(-701,32); cos_data_int <= to_signed(-713,32);
				when 2555 => sin_data_int <= to_signed(-702,32); cos_data_int <= to_signed(-711,32);
				when 2556 => sin_data_int <= to_signed(-703,32); cos_data_int <= to_signed(-710,32);
				when 2557 => sin_data_int <= to_signed(-704,32); cos_data_int <= to_signed(-709,32);
				when 2558 => sin_data_int <= to_signed(-705,32); cos_data_int <= to_signed(-708,32);
				when 2559 => sin_data_int <= to_signed(-706,32); cos_data_int <= to_signed(-707,32);
				when 2560 => sin_data_int <= to_signed(-707,32); cos_data_int <= to_signed(-706,32);
				when 2561 => sin_data_int <= to_signed(-708,32); cos_data_int <= to_signed(-705,32);
				when 2562 => sin_data_int <= to_signed(-709,32); cos_data_int <= to_signed(-704,32);
				when 2563 => sin_data_int <= to_signed(-710,32); cos_data_int <= to_signed(-703,32);
				when 2564 => sin_data_int <= to_signed(-711,32); cos_data_int <= to_signed(-702,32);
				when 2565 => sin_data_int <= to_signed(-713,32); cos_data_int <= to_signed(-701,32);
				when 2566 => sin_data_int <= to_signed(-714,32); cos_data_int <= to_signed(-699,32);
				when 2567 => sin_data_int <= to_signed(-715,32); cos_data_int <= to_signed(-698,32);
				when 2568 => sin_data_int <= to_signed(-716,32); cos_data_int <= to_signed(-697,32);
				when 2569 => sin_data_int <= to_signed(-717,32); cos_data_int <= to_signed(-696,32);
				when 2570 => sin_data_int <= to_signed(-718,32); cos_data_int <= to_signed(-695,32);
				when 2571 => sin_data_int <= to_signed(-719,32); cos_data_int <= to_signed(-694,32);
				when 2572 => sin_data_int <= to_signed(-720,32); cos_data_int <= to_signed(-693,32);
				when 2573 => sin_data_int <= to_signed(-721,32); cos_data_int <= to_signed(-692,32);
				when 2574 => sin_data_int <= to_signed(-722,32); cos_data_int <= to_signed(-691,32);
				when 2575 => sin_data_int <= to_signed(-723,32); cos_data_int <= to_signed(-690,32);
				when 2576 => sin_data_int <= to_signed(-724,32); cos_data_int <= to_signed(-688,32);
				when 2577 => sin_data_int <= to_signed(-725,32); cos_data_int <= to_signed(-687,32);
				when 2578 => sin_data_int <= to_signed(-726,32); cos_data_int <= to_signed(-686,32);
				when 2579 => sin_data_int <= to_signed(-727,32); cos_data_int <= to_signed(-685,32);
				when 2580 => sin_data_int <= to_signed(-728,32); cos_data_int <= to_signed(-684,32);
				when 2581 => sin_data_int <= to_signed(-730,32); cos_data_int <= to_signed(-683,32);
				when 2582 => sin_data_int <= to_signed(-731,32); cos_data_int <= to_signed(-682,32);
				when 2583 => sin_data_int <= to_signed(-732,32); cos_data_int <= to_signed(-681,32);
				when 2584 => sin_data_int <= to_signed(-733,32); cos_data_int <= to_signed(-679,32);
				when 2585 => sin_data_int <= to_signed(-734,32); cos_data_int <= to_signed(-678,32);
				when 2586 => sin_data_int <= to_signed(-735,32); cos_data_int <= to_signed(-677,32);
				when 2587 => sin_data_int <= to_signed(-736,32); cos_data_int <= to_signed(-676,32);
				when 2588 => sin_data_int <= to_signed(-737,32); cos_data_int <= to_signed(-675,32);
				when 2589 => sin_data_int <= to_signed(-738,32); cos_data_int <= to_signed(-674,32);
				when 2590 => sin_data_int <= to_signed(-739,32); cos_data_int <= to_signed(-673,32);
				when 2591 => sin_data_int <= to_signed(-740,32); cos_data_int <= to_signed(-672,32);
				when 2592 => sin_data_int <= to_signed(-741,32); cos_data_int <= to_signed(-670,32);
				when 2593 => sin_data_int <= to_signed(-742,32); cos_data_int <= to_signed(-669,32);
				when 2594 => sin_data_int <= to_signed(-743,32); cos_data_int <= to_signed(-668,32);
				when 2595 => sin_data_int <= to_signed(-744,32); cos_data_int <= to_signed(-667,32);
				when 2596 => sin_data_int <= to_signed(-745,32); cos_data_int <= to_signed(-666,32);
				when 2597 => sin_data_int <= to_signed(-746,32); cos_data_int <= to_signed(-665,32);
				when 2598 => sin_data_int <= to_signed(-747,32); cos_data_int <= to_signed(-664,32);
				when 2599 => sin_data_int <= to_signed(-748,32); cos_data_int <= to_signed(-662,32);
				when 2600 => sin_data_int <= to_signed(-749,32); cos_data_int <= to_signed(-661,32);
				when 2601 => sin_data_int <= to_signed(-750,32); cos_data_int <= to_signed(-660,32);
				when 2602 => sin_data_int <= to_signed(-751,32); cos_data_int <= to_signed(-659,32);
				when 2603 => sin_data_int <= to_signed(-752,32); cos_data_int <= to_signed(-658,32);
				when 2604 => sin_data_int <= to_signed(-753,32); cos_data_int <= to_signed(-657,32);
				when 2605 => sin_data_int <= to_signed(-754,32); cos_data_int <= to_signed(-655,32);
				when 2606 => sin_data_int <= to_signed(-755,32); cos_data_int <= to_signed(-654,32);
				when 2607 => sin_data_int <= to_signed(-756,32); cos_data_int <= to_signed(-653,32);
				when 2608 => sin_data_int <= to_signed(-757,32); cos_data_int <= to_signed(-652,32);
				when 2609 => sin_data_int <= to_signed(-758,32); cos_data_int <= to_signed(-651,32);
				when 2610 => sin_data_int <= to_signed(-759,32); cos_data_int <= to_signed(-650,32);
				when 2611 => sin_data_int <= to_signed(-760,32); cos_data_int <= to_signed(-649,32);
				when 2612 => sin_data_int <= to_signed(-761,32); cos_data_int <= to_signed(-647,32);
				when 2613 => sin_data_int <= to_signed(-762,32); cos_data_int <= to_signed(-646,32);
				when 2614 => sin_data_int <= to_signed(-763,32); cos_data_int <= to_signed(-645,32);
				when 2615 => sin_data_int <= to_signed(-764,32); cos_data_int <= to_signed(-644,32);
				when 2616 => sin_data_int <= to_signed(-765,32); cos_data_int <= to_signed(-643,32);
				when 2617 => sin_data_int <= to_signed(-766,32); cos_data_int <= to_signed(-641,32);
				when 2618 => sin_data_int <= to_signed(-767,32); cos_data_int <= to_signed(-640,32);
				when 2619 => sin_data_int <= to_signed(-768,32); cos_data_int <= to_signed(-639,32);
				when 2620 => sin_data_int <= to_signed(-769,32); cos_data_int <= to_signed(-638,32);
				when 2621 => sin_data_int <= to_signed(-770,32); cos_data_int <= to_signed(-637,32);
				when 2622 => sin_data_int <= to_signed(-771,32); cos_data_int <= to_signed(-636,32);
				when 2623 => sin_data_int <= to_signed(-772,32); cos_data_int <= to_signed(-634,32);
				when 2624 => sin_data_int <= to_signed(-773,32); cos_data_int <= to_signed(-633,32);
				when 2625 => sin_data_int <= to_signed(-774,32); cos_data_int <= to_signed(-632,32);
				when 2626 => sin_data_int <= to_signed(-775,32); cos_data_int <= to_signed(-631,32);
				when 2627 => sin_data_int <= to_signed(-776,32); cos_data_int <= to_signed(-630,32);
				when 2628 => sin_data_int <= to_signed(-777,32); cos_data_int <= to_signed(-628,32);
				when 2629 => sin_data_int <= to_signed(-778,32); cos_data_int <= to_signed(-627,32);
				when 2630 => sin_data_int <= to_signed(-779,32); cos_data_int <= to_signed(-626,32);
				when 2631 => sin_data_int <= to_signed(-780,32); cos_data_int <= to_signed(-625,32);
				when 2632 => sin_data_int <= to_signed(-781,32); cos_data_int <= to_signed(-624,32);
				when 2633 => sin_data_int <= to_signed(-782,32); cos_data_int <= to_signed(-622,32);
				when 2634 => sin_data_int <= to_signed(-783,32); cos_data_int <= to_signed(-621,32);
				when 2635 => sin_data_int <= to_signed(-784,32); cos_data_int <= to_signed(-620,32);
				when 2636 => sin_data_int <= to_signed(-785,32); cos_data_int <= to_signed(-619,32);
				when 2637 => sin_data_int <= to_signed(-786,32); cos_data_int <= to_signed(-618,32);
				when 2638 => sin_data_int <= to_signed(-786,32); cos_data_int <= to_signed(-616,32);
				when 2639 => sin_data_int <= to_signed(-787,32); cos_data_int <= to_signed(-615,32);
				when 2640 => sin_data_int <= to_signed(-788,32); cos_data_int <= to_signed(-614,32);
				when 2641 => sin_data_int <= to_signed(-789,32); cos_data_int <= to_signed(-613,32);
				when 2642 => sin_data_int <= to_signed(-790,32); cos_data_int <= to_signed(-612,32);
				when 2643 => sin_data_int <= to_signed(-791,32); cos_data_int <= to_signed(-610,32);
				when 2644 => sin_data_int <= to_signed(-792,32); cos_data_int <= to_signed(-609,32);
				when 2645 => sin_data_int <= to_signed(-793,32); cos_data_int <= to_signed(-608,32);
				when 2646 => sin_data_int <= to_signed(-794,32); cos_data_int <= to_signed(-607,32);
				when 2647 => sin_data_int <= to_signed(-795,32); cos_data_int <= to_signed(-606,32);
				when 2648 => sin_data_int <= to_signed(-796,32); cos_data_int <= to_signed(-604,32);
				when 2649 => sin_data_int <= to_signed(-797,32); cos_data_int <= to_signed(-603,32);
				when 2650 => sin_data_int <= to_signed(-798,32); cos_data_int <= to_signed(-602,32);
				when 2651 => sin_data_int <= to_signed(-799,32); cos_data_int <= to_signed(-601,32);
				when 2652 => sin_data_int <= to_signed(-800,32); cos_data_int <= to_signed(-599,32);
				when 2653 => sin_data_int <= to_signed(-800,32); cos_data_int <= to_signed(-598,32);
				when 2654 => sin_data_int <= to_signed(-801,32); cos_data_int <= to_signed(-597,32);
				when 2655 => sin_data_int <= to_signed(-802,32); cos_data_int <= to_signed(-596,32);
				when 2656 => sin_data_int <= to_signed(-803,32); cos_data_int <= to_signed(-594,32);
				when 2657 => sin_data_int <= to_signed(-804,32); cos_data_int <= to_signed(-593,32);
				when 2658 => sin_data_int <= to_signed(-805,32); cos_data_int <= to_signed(-592,32);
				when 2659 => sin_data_int <= to_signed(-806,32); cos_data_int <= to_signed(-591,32);
				when 2660 => sin_data_int <= to_signed(-807,32); cos_data_int <= to_signed(-590,32);
				when 2661 => sin_data_int <= to_signed(-808,32); cos_data_int <= to_signed(-588,32);
				when 2662 => sin_data_int <= to_signed(-809,32); cos_data_int <= to_signed(-587,32);
				when 2663 => sin_data_int <= to_signed(-810,32); cos_data_int <= to_signed(-586,32);
				when 2664 => sin_data_int <= to_signed(-810,32); cos_data_int <= to_signed(-585,32);
				when 2665 => sin_data_int <= to_signed(-811,32); cos_data_int <= to_signed(-583,32);
				when 2666 => sin_data_int <= to_signed(-812,32); cos_data_int <= to_signed(-582,32);
				when 2667 => sin_data_int <= to_signed(-813,32); cos_data_int <= to_signed(-581,32);
				when 2668 => sin_data_int <= to_signed(-814,32); cos_data_int <= to_signed(-580,32);
				when 2669 => sin_data_int <= to_signed(-815,32); cos_data_int <= to_signed(-578,32);
				when 2670 => sin_data_int <= to_signed(-816,32); cos_data_int <= to_signed(-577,32);
				when 2671 => sin_data_int <= to_signed(-817,32); cos_data_int <= to_signed(-576,32);
				when 2672 => sin_data_int <= to_signed(-818,32); cos_data_int <= to_signed(-575,32);
				when 2673 => sin_data_int <= to_signed(-818,32); cos_data_int <= to_signed(-573,32);
				when 2674 => sin_data_int <= to_signed(-819,32); cos_data_int <= to_signed(-572,32);
				when 2675 => sin_data_int <= to_signed(-820,32); cos_data_int <= to_signed(-571,32);
				when 2676 => sin_data_int <= to_signed(-821,32); cos_data_int <= to_signed(-570,32);
				when 2677 => sin_data_int <= to_signed(-822,32); cos_data_int <= to_signed(-568,32);
				when 2678 => sin_data_int <= to_signed(-823,32); cos_data_int <= to_signed(-567,32);
				when 2679 => sin_data_int <= to_signed(-824,32); cos_data_int <= to_signed(-566,32);
				when 2680 => sin_data_int <= to_signed(-825,32); cos_data_int <= to_signed(-564,32);
				when 2681 => sin_data_int <= to_signed(-825,32); cos_data_int <= to_signed(-563,32);
				when 2682 => sin_data_int <= to_signed(-826,32); cos_data_int <= to_signed(-562,32);
				when 2683 => sin_data_int <= to_signed(-827,32); cos_data_int <= to_signed(-561,32);
				when 2684 => sin_data_int <= to_signed(-828,32); cos_data_int <= to_signed(-559,32);
				when 2685 => sin_data_int <= to_signed(-829,32); cos_data_int <= to_signed(-558,32);
				when 2686 => sin_data_int <= to_signed(-830,32); cos_data_int <= to_signed(-557,32);
				when 2687 => sin_data_int <= to_signed(-831,32); cos_data_int <= to_signed(-556,32);
				when 2688 => sin_data_int <= to_signed(-831,32); cos_data_int <= to_signed(-554,32);
				when 2689 => sin_data_int <= to_signed(-832,32); cos_data_int <= to_signed(-553,32);
				when 2690 => sin_data_int <= to_signed(-833,32); cos_data_int <= to_signed(-552,32);
				when 2691 => sin_data_int <= to_signed(-834,32); cos_data_int <= to_signed(-550,32);
				when 2692 => sin_data_int <= to_signed(-835,32); cos_data_int <= to_signed(-549,32);
				when 2693 => sin_data_int <= to_signed(-836,32); cos_data_int <= to_signed(-548,32);
				when 2694 => sin_data_int <= to_signed(-837,32); cos_data_int <= to_signed(-547,32);
				when 2695 => sin_data_int <= to_signed(-837,32); cos_data_int <= to_signed(-545,32);
				when 2696 => sin_data_int <= to_signed(-838,32); cos_data_int <= to_signed(-544,32);
				when 2697 => sin_data_int <= to_signed(-839,32); cos_data_int <= to_signed(-543,32);
				when 2698 => sin_data_int <= to_signed(-840,32); cos_data_int <= to_signed(-541,32);
				when 2699 => sin_data_int <= to_signed(-841,32); cos_data_int <= to_signed(-540,32);
				when 2700 => sin_data_int <= to_signed(-842,32); cos_data_int <= to_signed(-539,32);
				when 2701 => sin_data_int <= to_signed(-842,32); cos_data_int <= to_signed(-538,32);
				when 2702 => sin_data_int <= to_signed(-843,32); cos_data_int <= to_signed(-536,32);
				when 2703 => sin_data_int <= to_signed(-844,32); cos_data_int <= to_signed(-535,32);
				when 2704 => sin_data_int <= to_signed(-845,32); cos_data_int <= to_signed(-534,32);
				when 2705 => sin_data_int <= to_signed(-846,32); cos_data_int <= to_signed(-532,32);
				when 2706 => sin_data_int <= to_signed(-846,32); cos_data_int <= to_signed(-531,32);
				when 2707 => sin_data_int <= to_signed(-847,32); cos_data_int <= to_signed(-530,32);
				when 2708 => sin_data_int <= to_signed(-848,32); cos_data_int <= to_signed(-529,32);
				when 2709 => sin_data_int <= to_signed(-849,32); cos_data_int <= to_signed(-527,32);
				when 2710 => sin_data_int <= to_signed(-850,32); cos_data_int <= to_signed(-526,32);
				when 2711 => sin_data_int <= to_signed(-851,32); cos_data_int <= to_signed(-525,32);
				when 2712 => sin_data_int <= to_signed(-851,32); cos_data_int <= to_signed(-523,32);
				when 2713 => sin_data_int <= to_signed(-852,32); cos_data_int <= to_signed(-522,32);
				when 2714 => sin_data_int <= to_signed(-853,32); cos_data_int <= to_signed(-521,32);
				when 2715 => sin_data_int <= to_signed(-854,32); cos_data_int <= to_signed(-519,32);
				when 2716 => sin_data_int <= to_signed(-855,32); cos_data_int <= to_signed(-518,32);
				when 2717 => sin_data_int <= to_signed(-855,32); cos_data_int <= to_signed(-517,32);
				when 2718 => sin_data_int <= to_signed(-856,32); cos_data_int <= to_signed(-515,32);
				when 2719 => sin_data_int <= to_signed(-857,32); cos_data_int <= to_signed(-514,32);
				when 2720 => sin_data_int <= to_signed(-858,32); cos_data_int <= to_signed(-513,32);
				when 2721 => sin_data_int <= to_signed(-859,32); cos_data_int <= to_signed(-511,32);
				when 2722 => sin_data_int <= to_signed(-859,32); cos_data_int <= to_signed(-510,32);
				when 2723 => sin_data_int <= to_signed(-860,32); cos_data_int <= to_signed(-509,32);
				when 2724 => sin_data_int <= to_signed(-861,32); cos_data_int <= to_signed(-508,32);
				when 2725 => sin_data_int <= to_signed(-862,32); cos_data_int <= to_signed(-506,32);
				when 2726 => sin_data_int <= to_signed(-862,32); cos_data_int <= to_signed(-505,32);
				when 2727 => sin_data_int <= to_signed(-863,32); cos_data_int <= to_signed(-504,32);
				when 2728 => sin_data_int <= to_signed(-864,32); cos_data_int <= to_signed(-502,32);
				when 2729 => sin_data_int <= to_signed(-865,32); cos_data_int <= to_signed(-501,32);
				when 2730 => sin_data_int <= to_signed(-866,32); cos_data_int <= to_signed(-500,32);
				when 2731 => sin_data_int <= to_signed(-866,32); cos_data_int <= to_signed(-498,32);
				when 2732 => sin_data_int <= to_signed(-867,32); cos_data_int <= to_signed(-497,32);
				when 2733 => sin_data_int <= to_signed(-868,32); cos_data_int <= to_signed(-496,32);
				when 2734 => sin_data_int <= to_signed(-869,32); cos_data_int <= to_signed(-494,32);
				when 2735 => sin_data_int <= to_signed(-869,32); cos_data_int <= to_signed(-493,32);
				when 2736 => sin_data_int <= to_signed(-870,32); cos_data_int <= to_signed(-492,32);
				when 2737 => sin_data_int <= to_signed(-871,32); cos_data_int <= to_signed(-490,32);
				when 2738 => sin_data_int <= to_signed(-872,32); cos_data_int <= to_signed(-489,32);
				when 2739 => sin_data_int <= to_signed(-872,32); cos_data_int <= to_signed(-488,32);
				when 2740 => sin_data_int <= to_signed(-873,32); cos_data_int <= to_signed(-486,32);
				when 2741 => sin_data_int <= to_signed(-874,32); cos_data_int <= to_signed(-485,32);
				when 2742 => sin_data_int <= to_signed(-875,32); cos_data_int <= to_signed(-484,32);
				when 2743 => sin_data_int <= to_signed(-875,32); cos_data_int <= to_signed(-482,32);
				when 2744 => sin_data_int <= to_signed(-876,32); cos_data_int <= to_signed(-481,32);
				when 2745 => sin_data_int <= to_signed(-877,32); cos_data_int <= to_signed(-479,32);
				when 2746 => sin_data_int <= to_signed(-878,32); cos_data_int <= to_signed(-478,32);
				when 2747 => sin_data_int <= to_signed(-878,32); cos_data_int <= to_signed(-477,32);
				when 2748 => sin_data_int <= to_signed(-879,32); cos_data_int <= to_signed(-475,32);
				when 2749 => sin_data_int <= to_signed(-880,32); cos_data_int <= to_signed(-474,32);
				when 2750 => sin_data_int <= to_signed(-880,32); cos_data_int <= to_signed(-473,32);
				when 2751 => sin_data_int <= to_signed(-881,32); cos_data_int <= to_signed(-471,32);
				when 2752 => sin_data_int <= to_signed(-882,32); cos_data_int <= to_signed(-470,32);
				when 2753 => sin_data_int <= to_signed(-883,32); cos_data_int <= to_signed(-469,32);
				when 2754 => sin_data_int <= to_signed(-883,32); cos_data_int <= to_signed(-467,32);
				when 2755 => sin_data_int <= to_signed(-884,32); cos_data_int <= to_signed(-466,32);
				when 2756 => sin_data_int <= to_signed(-885,32); cos_data_int <= to_signed(-465,32);
				when 2757 => sin_data_int <= to_signed(-886,32); cos_data_int <= to_signed(-463,32);
				when 2758 => sin_data_int <= to_signed(-886,32); cos_data_int <= to_signed(-462,32);
				when 2759 => sin_data_int <= to_signed(-887,32); cos_data_int <= to_signed(-461,32);
				when 2760 => sin_data_int <= to_signed(-888,32); cos_data_int <= to_signed(-459,32);
				when 2761 => sin_data_int <= to_signed(-888,32); cos_data_int <= to_signed(-458,32);
				when 2762 => sin_data_int <= to_signed(-889,32); cos_data_int <= to_signed(-456,32);
				when 2763 => sin_data_int <= to_signed(-890,32); cos_data_int <= to_signed(-455,32);
				when 2764 => sin_data_int <= to_signed(-890,32); cos_data_int <= to_signed(-454,32);
				when 2765 => sin_data_int <= to_signed(-891,32); cos_data_int <= to_signed(-452,32);
				when 2766 => sin_data_int <= to_signed(-892,32); cos_data_int <= to_signed(-451,32);
				when 2767 => sin_data_int <= to_signed(-893,32); cos_data_int <= to_signed(-450,32);
				when 2768 => sin_data_int <= to_signed(-893,32); cos_data_int <= to_signed(-448,32);
				when 2769 => sin_data_int <= to_signed(-894,32); cos_data_int <= to_signed(-447,32);
				when 2770 => sin_data_int <= to_signed(-895,32); cos_data_int <= to_signed(-445,32);
				when 2771 => sin_data_int <= to_signed(-895,32); cos_data_int <= to_signed(-444,32);
				when 2772 => sin_data_int <= to_signed(-896,32); cos_data_int <= to_signed(-443,32);
				when 2773 => sin_data_int <= to_signed(-897,32); cos_data_int <= to_signed(-441,32);
				when 2774 => sin_data_int <= to_signed(-897,32); cos_data_int <= to_signed(-440,32);
				when 2775 => sin_data_int <= to_signed(-898,32); cos_data_int <= to_signed(-439,32);
				when 2776 => sin_data_int <= to_signed(-899,32); cos_data_int <= to_signed(-437,32);
				when 2777 => sin_data_int <= to_signed(-899,32); cos_data_int <= to_signed(-436,32);
				when 2778 => sin_data_int <= to_signed(-900,32); cos_data_int <= to_signed(-434,32);
				when 2779 => sin_data_int <= to_signed(-901,32); cos_data_int <= to_signed(-433,32);
				when 2780 => sin_data_int <= to_signed(-901,32); cos_data_int <= to_signed(-432,32);
				when 2781 => sin_data_int <= to_signed(-902,32); cos_data_int <= to_signed(-430,32);
				when 2782 => sin_data_int <= to_signed(-903,32); cos_data_int <= to_signed(-429,32);
				when 2783 => sin_data_int <= to_signed(-903,32); cos_data_int <= to_signed(-428,32);
				when 2784 => sin_data_int <= to_signed(-904,32); cos_data_int <= to_signed(-426,32);
				when 2785 => sin_data_int <= to_signed(-905,32); cos_data_int <= to_signed(-425,32);
				when 2786 => sin_data_int <= to_signed(-905,32); cos_data_int <= to_signed(-423,32);
				when 2787 => sin_data_int <= to_signed(-906,32); cos_data_int <= to_signed(-422,32);
				when 2788 => sin_data_int <= to_signed(-907,32); cos_data_int <= to_signed(-421,32);
				when 2789 => sin_data_int <= to_signed(-907,32); cos_data_int <= to_signed(-419,32);
				when 2790 => sin_data_int <= to_signed(-908,32); cos_data_int <= to_signed(-418,32);
				when 2791 => sin_data_int <= to_signed(-909,32); cos_data_int <= to_signed(-416,32);
				when 2792 => sin_data_int <= to_signed(-909,32); cos_data_int <= to_signed(-415,32);
				when 2793 => sin_data_int <= to_signed(-910,32); cos_data_int <= to_signed(-414,32);
				when 2794 => sin_data_int <= to_signed(-910,32); cos_data_int <= to_signed(-412,32);
				when 2795 => sin_data_int <= to_signed(-911,32); cos_data_int <= to_signed(-411,32);
				when 2796 => sin_data_int <= to_signed(-912,32); cos_data_int <= to_signed(-409,32);
				when 2797 => sin_data_int <= to_signed(-912,32); cos_data_int <= to_signed(-408,32);
				when 2798 => sin_data_int <= to_signed(-913,32); cos_data_int <= to_signed(-407,32);
				when 2799 => sin_data_int <= to_signed(-914,32); cos_data_int <= to_signed(-405,32);
				when 2800 => sin_data_int <= to_signed(-914,32); cos_data_int <= to_signed(-404,32);
				when 2801 => sin_data_int <= to_signed(-915,32); cos_data_int <= to_signed(-402,32);
				when 2802 => sin_data_int <= to_signed(-915,32); cos_data_int <= to_signed(-401,32);
				when 2803 => sin_data_int <= to_signed(-916,32); cos_data_int <= to_signed(-400,32);
				when 2804 => sin_data_int <= to_signed(-917,32); cos_data_int <= to_signed(-398,32);
				when 2805 => sin_data_int <= to_signed(-917,32); cos_data_int <= to_signed(-397,32);
				when 2806 => sin_data_int <= to_signed(-918,32); cos_data_int <= to_signed(-395,32);
				when 2807 => sin_data_int <= to_signed(-919,32); cos_data_int <= to_signed(-394,32);
				when 2808 => sin_data_int <= to_signed(-919,32); cos_data_int <= to_signed(-393,32);
				when 2809 => sin_data_int <= to_signed(-920,32); cos_data_int <= to_signed(-391,32);
				when 2810 => sin_data_int <= to_signed(-920,32); cos_data_int <= to_signed(-390,32);
				when 2811 => sin_data_int <= to_signed(-921,32); cos_data_int <= to_signed(-388,32);
				when 2812 => sin_data_int <= to_signed(-922,32); cos_data_int <= to_signed(-387,32);
				when 2813 => sin_data_int <= to_signed(-922,32); cos_data_int <= to_signed(-386,32);
				when 2814 => sin_data_int <= to_signed(-923,32); cos_data_int <= to_signed(-384,32);
				when 2815 => sin_data_int <= to_signed(-923,32); cos_data_int <= to_signed(-383,32);
				when 2816 => sin_data_int <= to_signed(-924,32); cos_data_int <= to_signed(-381,32);
				when 2817 => sin_data_int <= to_signed(-924,32); cos_data_int <= to_signed(-380,32);
				when 2818 => sin_data_int <= to_signed(-925,32); cos_data_int <= to_signed(-378,32);
				when 2819 => sin_data_int <= to_signed(-926,32); cos_data_int <= to_signed(-377,32);
				when 2820 => sin_data_int <= to_signed(-926,32); cos_data_int <= to_signed(-376,32);
				when 2821 => sin_data_int <= to_signed(-927,32); cos_data_int <= to_signed(-374,32);
				when 2822 => sin_data_int <= to_signed(-927,32); cos_data_int <= to_signed(-373,32);
				when 2823 => sin_data_int <= to_signed(-928,32); cos_data_int <= to_signed(-371,32);
				when 2824 => sin_data_int <= to_signed(-929,32); cos_data_int <= to_signed(-370,32);
				when 2825 => sin_data_int <= to_signed(-929,32); cos_data_int <= to_signed(-368,32);
				when 2826 => sin_data_int <= to_signed(-930,32); cos_data_int <= to_signed(-367,32);
				when 2827 => sin_data_int <= to_signed(-930,32); cos_data_int <= to_signed(-366,32);
				when 2828 => sin_data_int <= to_signed(-931,32); cos_data_int <= to_signed(-364,32);
				when 2829 => sin_data_int <= to_signed(-931,32); cos_data_int <= to_signed(-363,32);
				when 2830 => sin_data_int <= to_signed(-932,32); cos_data_int <= to_signed(-361,32);
				when 2831 => sin_data_int <= to_signed(-932,32); cos_data_int <= to_signed(-360,32);
				when 2832 => sin_data_int <= to_signed(-933,32); cos_data_int <= to_signed(-358,32);
				when 2833 => sin_data_int <= to_signed(-934,32); cos_data_int <= to_signed(-357,32);
				when 2834 => sin_data_int <= to_signed(-934,32); cos_data_int <= to_signed(-356,32);
				when 2835 => sin_data_int <= to_signed(-935,32); cos_data_int <= to_signed(-354,32);
				when 2836 => sin_data_int <= to_signed(-935,32); cos_data_int <= to_signed(-353,32);
				when 2837 => sin_data_int <= to_signed(-936,32); cos_data_int <= to_signed(-351,32);
				when 2838 => sin_data_int <= to_signed(-936,32); cos_data_int <= to_signed(-350,32);
				when 2839 => sin_data_int <= to_signed(-937,32); cos_data_int <= to_signed(-348,32);
				when 2840 => sin_data_int <= to_signed(-937,32); cos_data_int <= to_signed(-347,32);
				when 2841 => sin_data_int <= to_signed(-938,32); cos_data_int <= to_signed(-346,32);
				when 2842 => sin_data_int <= to_signed(-938,32); cos_data_int <= to_signed(-344,32);
				when 2843 => sin_data_int <= to_signed(-939,32); cos_data_int <= to_signed(-343,32);
				when 2844 => sin_data_int <= to_signed(-939,32); cos_data_int <= to_signed(-341,32);
				when 2845 => sin_data_int <= to_signed(-940,32); cos_data_int <= to_signed(-340,32);
				when 2846 => sin_data_int <= to_signed(-941,32); cos_data_int <= to_signed(-338,32);
				when 2847 => sin_data_int <= to_signed(-941,32); cos_data_int <= to_signed(-337,32);
				when 2848 => sin_data_int <= to_signed(-942,32); cos_data_int <= to_signed(-335,32);
				when 2849 => sin_data_int <= to_signed(-942,32); cos_data_int <= to_signed(-334,32);
				when 2850 => sin_data_int <= to_signed(-943,32); cos_data_int <= to_signed(-333,32);
				when 2851 => sin_data_int <= to_signed(-943,32); cos_data_int <= to_signed(-331,32);
				when 2852 => sin_data_int <= to_signed(-944,32); cos_data_int <= to_signed(-330,32);
				when 2853 => sin_data_int <= to_signed(-944,32); cos_data_int <= to_signed(-328,32);
				when 2854 => sin_data_int <= to_signed(-945,32); cos_data_int <= to_signed(-327,32);
				when 2855 => sin_data_int <= to_signed(-945,32); cos_data_int <= to_signed(-325,32);
				when 2856 => sin_data_int <= to_signed(-946,32); cos_data_int <= to_signed(-324,32);
				when 2857 => sin_data_int <= to_signed(-946,32); cos_data_int <= to_signed(-322,32);
				when 2858 => sin_data_int <= to_signed(-947,32); cos_data_int <= to_signed(-321,32);
				when 2859 => sin_data_int <= to_signed(-947,32); cos_data_int <= to_signed(-320,32);
				when 2860 => sin_data_int <= to_signed(-948,32); cos_data_int <= to_signed(-318,32);
				when 2861 => sin_data_int <= to_signed(-948,32); cos_data_int <= to_signed(-317,32);
				when 2862 => sin_data_int <= to_signed(-949,32); cos_data_int <= to_signed(-315,32);
				when 2863 => sin_data_int <= to_signed(-949,32); cos_data_int <= to_signed(-314,32);
				when 2864 => sin_data_int <= to_signed(-950,32); cos_data_int <= to_signed(-312,32);
				when 2865 => sin_data_int <= to_signed(-950,32); cos_data_int <= to_signed(-311,32);
				when 2866 => sin_data_int <= to_signed(-950,32); cos_data_int <= to_signed(-309,32);
				when 2867 => sin_data_int <= to_signed(-951,32); cos_data_int <= to_signed(-308,32);
				when 2868 => sin_data_int <= to_signed(-951,32); cos_data_int <= to_signed(-306,32);
				when 2869 => sin_data_int <= to_signed(-952,32); cos_data_int <= to_signed(-305,32);
				when 2870 => sin_data_int <= to_signed(-952,32); cos_data_int <= to_signed(-303,32);
				when 2871 => sin_data_int <= to_signed(-953,32); cos_data_int <= to_signed(-302,32);
				when 2872 => sin_data_int <= to_signed(-953,32); cos_data_int <= to_signed(-301,32);
				when 2873 => sin_data_int <= to_signed(-954,32); cos_data_int <= to_signed(-299,32);
				when 2874 => sin_data_int <= to_signed(-954,32); cos_data_int <= to_signed(-298,32);
				when 2875 => sin_data_int <= to_signed(-955,32); cos_data_int <= to_signed(-296,32);
				when 2876 => sin_data_int <= to_signed(-955,32); cos_data_int <= to_signed(-295,32);
				when 2877 => sin_data_int <= to_signed(-956,32); cos_data_int <= to_signed(-293,32);
				when 2878 => sin_data_int <= to_signed(-956,32); cos_data_int <= to_signed(-292,32);
				when 2879 => sin_data_int <= to_signed(-956,32); cos_data_int <= to_signed(-290,32);
				when 2880 => sin_data_int <= to_signed(-957,32); cos_data_int <= to_signed(-289,32);
				when 2881 => sin_data_int <= to_signed(-957,32); cos_data_int <= to_signed(-287,32);
				when 2882 => sin_data_int <= to_signed(-958,32); cos_data_int <= to_signed(-286,32);
				when 2883 => sin_data_int <= to_signed(-958,32); cos_data_int <= to_signed(-284,32);
				when 2884 => sin_data_int <= to_signed(-959,32); cos_data_int <= to_signed(-283,32);
				when 2885 => sin_data_int <= to_signed(-959,32); cos_data_int <= to_signed(-281,32);
				when 2886 => sin_data_int <= to_signed(-960,32); cos_data_int <= to_signed(-280,32);
				when 2887 => sin_data_int <= to_signed(-960,32); cos_data_int <= to_signed(-279,32);
				when 2888 => sin_data_int <= to_signed(-960,32); cos_data_int <= to_signed(-277,32);
				when 2889 => sin_data_int <= to_signed(-961,32); cos_data_int <= to_signed(-276,32);
				when 2890 => sin_data_int <= to_signed(-961,32); cos_data_int <= to_signed(-274,32);
				when 2891 => sin_data_int <= to_signed(-962,32); cos_data_int <= to_signed(-273,32);
				when 2892 => sin_data_int <= to_signed(-962,32); cos_data_int <= to_signed(-271,32);
				when 2893 => sin_data_int <= to_signed(-963,32); cos_data_int <= to_signed(-270,32);
				when 2894 => sin_data_int <= to_signed(-963,32); cos_data_int <= to_signed(-268,32);
				when 2895 => sin_data_int <= to_signed(-963,32); cos_data_int <= to_signed(-267,32);
				when 2896 => sin_data_int <= to_signed(-964,32); cos_data_int <= to_signed(-265,32);
				when 2897 => sin_data_int <= to_signed(-964,32); cos_data_int <= to_signed(-264,32);
				when 2898 => sin_data_int <= to_signed(-965,32); cos_data_int <= to_signed(-262,32);
				when 2899 => sin_data_int <= to_signed(-965,32); cos_data_int <= to_signed(-261,32);
				when 2900 => sin_data_int <= to_signed(-965,32); cos_data_int <= to_signed(-259,32);
				when 2901 => sin_data_int <= to_signed(-966,32); cos_data_int <= to_signed(-258,32);
				when 2902 => sin_data_int <= to_signed(-966,32); cos_data_int <= to_signed(-256,32);
				when 2903 => sin_data_int <= to_signed(-967,32); cos_data_int <= to_signed(-255,32);
				when 2904 => sin_data_int <= to_signed(-967,32); cos_data_int <= to_signed(-253,32);
				when 2905 => sin_data_int <= to_signed(-967,32); cos_data_int <= to_signed(-252,32);
				when 2906 => sin_data_int <= to_signed(-968,32); cos_data_int <= to_signed(-250,32);
				when 2907 => sin_data_int <= to_signed(-968,32); cos_data_int <= to_signed(-249,32);
				when 2908 => sin_data_int <= to_signed(-969,32); cos_data_int <= to_signed(-247,32);
				when 2909 => sin_data_int <= to_signed(-969,32); cos_data_int <= to_signed(-246,32);
				when 2910 => sin_data_int <= to_signed(-969,32); cos_data_int <= to_signed(-244,32);
				when 2911 => sin_data_int <= to_signed(-970,32); cos_data_int <= to_signed(-243,32);
				when 2912 => sin_data_int <= to_signed(-970,32); cos_data_int <= to_signed(-241,32);
				when 2913 => sin_data_int <= to_signed(-970,32); cos_data_int <= to_signed(-240,32);
				when 2914 => sin_data_int <= to_signed(-971,32); cos_data_int <= to_signed(-239,32);
				when 2915 => sin_data_int <= to_signed(-971,32); cos_data_int <= to_signed(-237,32);
				when 2916 => sin_data_int <= to_signed(-972,32); cos_data_int <= to_signed(-236,32);
				when 2917 => sin_data_int <= to_signed(-972,32); cos_data_int <= to_signed(-234,32);
				when 2918 => sin_data_int <= to_signed(-972,32); cos_data_int <= to_signed(-233,32);
				when 2919 => sin_data_int <= to_signed(-973,32); cos_data_int <= to_signed(-231,32);
				when 2920 => sin_data_int <= to_signed(-973,32); cos_data_int <= to_signed(-230,32);
				when 2921 => sin_data_int <= to_signed(-973,32); cos_data_int <= to_signed(-228,32);
				when 2922 => sin_data_int <= to_signed(-974,32); cos_data_int <= to_signed(-227,32);
				when 2923 => sin_data_int <= to_signed(-974,32); cos_data_int <= to_signed(-225,32);
				when 2924 => sin_data_int <= to_signed(-974,32); cos_data_int <= to_signed(-224,32);
				when 2925 => sin_data_int <= to_signed(-975,32); cos_data_int <= to_signed(-222,32);
				when 2926 => sin_data_int <= to_signed(-975,32); cos_data_int <= to_signed(-221,32);
				when 2927 => sin_data_int <= to_signed(-975,32); cos_data_int <= to_signed(-219,32);
				when 2928 => sin_data_int <= to_signed(-976,32); cos_data_int <= to_signed(-218,32);
				when 2929 => sin_data_int <= to_signed(-976,32); cos_data_int <= to_signed(-216,32);
				when 2930 => sin_data_int <= to_signed(-976,32); cos_data_int <= to_signed(-215,32);
				when 2931 => sin_data_int <= to_signed(-977,32); cos_data_int <= to_signed(-213,32);
				when 2932 => sin_data_int <= to_signed(-977,32); cos_data_int <= to_signed(-212,32);
				when 2933 => sin_data_int <= to_signed(-977,32); cos_data_int <= to_signed(-210,32);
				when 2934 => sin_data_int <= to_signed(-978,32); cos_data_int <= to_signed(-209,32);
				when 2935 => sin_data_int <= to_signed(-978,32); cos_data_int <= to_signed(-207,32);
				when 2936 => sin_data_int <= to_signed(-978,32); cos_data_int <= to_signed(-206,32);
				when 2937 => sin_data_int <= to_signed(-979,32); cos_data_int <= to_signed(-204,32);
				when 2938 => sin_data_int <= to_signed(-979,32); cos_data_int <= to_signed(-203,32);
				when 2939 => sin_data_int <= to_signed(-979,32); cos_data_int <= to_signed(-201,32);
				when 2940 => sin_data_int <= to_signed(-980,32); cos_data_int <= to_signed(-200,32);
				when 2941 => sin_data_int <= to_signed(-980,32); cos_data_int <= to_signed(-198,32);
				when 2942 => sin_data_int <= to_signed(-980,32); cos_data_int <= to_signed(-197,32);
				when 2943 => sin_data_int <= to_signed(-980,32); cos_data_int <= to_signed(-195,32);
				when 2944 => sin_data_int <= to_signed(-981,32); cos_data_int <= to_signed(-194,32);
				when 2945 => sin_data_int <= to_signed(-981,32); cos_data_int <= to_signed(-192,32);
				when 2946 => sin_data_int <= to_signed(-981,32); cos_data_int <= to_signed(-191,32);
				when 2947 => sin_data_int <= to_signed(-982,32); cos_data_int <= to_signed(-189,32);
				when 2948 => sin_data_int <= to_signed(-982,32); cos_data_int <= to_signed(-188,32);
				when 2949 => sin_data_int <= to_signed(-982,32); cos_data_int <= to_signed(-186,32);
				when 2950 => sin_data_int <= to_signed(-983,32); cos_data_int <= to_signed(-185,32);
				when 2951 => sin_data_int <= to_signed(-983,32); cos_data_int <= to_signed(-183,32);
				when 2952 => sin_data_int <= to_signed(-983,32); cos_data_int <= to_signed(-182,32);
				when 2953 => sin_data_int <= to_signed(-983,32); cos_data_int <= to_signed(-180,32);
				when 2954 => sin_data_int <= to_signed(-984,32); cos_data_int <= to_signed(-179,32);
				when 2955 => sin_data_int <= to_signed(-984,32); cos_data_int <= to_signed(-177,32);
				when 2956 => sin_data_int <= to_signed(-984,32); cos_data_int <= to_signed(-175,32);
				when 2957 => sin_data_int <= to_signed(-984,32); cos_data_int <= to_signed(-174,32);
				when 2958 => sin_data_int <= to_signed(-985,32); cos_data_int <= to_signed(-172,32);
				when 2959 => sin_data_int <= to_signed(-985,32); cos_data_int <= to_signed(-171,32);
				when 2960 => sin_data_int <= to_signed(-985,32); cos_data_int <= to_signed(-169,32);
				when 2961 => sin_data_int <= to_signed(-986,32); cos_data_int <= to_signed(-168,32);
				when 2962 => sin_data_int <= to_signed(-986,32); cos_data_int <= to_signed(-166,32);
				when 2963 => sin_data_int <= to_signed(-986,32); cos_data_int <= to_signed(-165,32);
				when 2964 => sin_data_int <= to_signed(-986,32); cos_data_int <= to_signed(-163,32);
				when 2965 => sin_data_int <= to_signed(-987,32); cos_data_int <= to_signed(-162,32);
				when 2966 => sin_data_int <= to_signed(-987,32); cos_data_int <= to_signed(-160,32);
				when 2967 => sin_data_int <= to_signed(-987,32); cos_data_int <= to_signed(-159,32);
				when 2968 => sin_data_int <= to_signed(-987,32); cos_data_int <= to_signed(-157,32);
				when 2969 => sin_data_int <= to_signed(-988,32); cos_data_int <= to_signed(-156,32);
				when 2970 => sin_data_int <= to_signed(-988,32); cos_data_int <= to_signed(-154,32);
				when 2971 => sin_data_int <= to_signed(-988,32); cos_data_int <= to_signed(-153,32);
				when 2972 => sin_data_int <= to_signed(-988,32); cos_data_int <= to_signed(-151,32);
				when 2973 => sin_data_int <= to_signed(-988,32); cos_data_int <= to_signed(-150,32);
				when 2974 => sin_data_int <= to_signed(-989,32); cos_data_int <= to_signed(-148,32);
				when 2975 => sin_data_int <= to_signed(-989,32); cos_data_int <= to_signed(-147,32);
				when 2976 => sin_data_int <= to_signed(-989,32); cos_data_int <= to_signed(-145,32);
				when 2977 => sin_data_int <= to_signed(-989,32); cos_data_int <= to_signed(-144,32);
				when 2978 => sin_data_int <= to_signed(-990,32); cos_data_int <= to_signed(-142,32);
				when 2979 => sin_data_int <= to_signed(-990,32); cos_data_int <= to_signed(-141,32);
				when 2980 => sin_data_int <= to_signed(-990,32); cos_data_int <= to_signed(-139,32);
				when 2981 => sin_data_int <= to_signed(-990,32); cos_data_int <= to_signed(-138,32);
				when 2982 => sin_data_int <= to_signed(-990,32); cos_data_int <= to_signed(-136,32);
				when 2983 => sin_data_int <= to_signed(-991,32); cos_data_int <= to_signed(-135,32);
				when 2984 => sin_data_int <= to_signed(-991,32); cos_data_int <= to_signed(-133,32);
				when 2985 => sin_data_int <= to_signed(-991,32); cos_data_int <= to_signed(-132,32);
				when 2986 => sin_data_int <= to_signed(-991,32); cos_data_int <= to_signed(-130,32);
				when 2987 => sin_data_int <= to_signed(-992,32); cos_data_int <= to_signed(-128,32);
				when 2988 => sin_data_int <= to_signed(-992,32); cos_data_int <= to_signed(-127,32);
				when 2989 => sin_data_int <= to_signed(-992,32); cos_data_int <= to_signed(-125,32);
				when 2990 => sin_data_int <= to_signed(-992,32); cos_data_int <= to_signed(-124,32);
				when 2991 => sin_data_int <= to_signed(-992,32); cos_data_int <= to_signed(-122,32);
				when 2992 => sin_data_int <= to_signed(-992,32); cos_data_int <= to_signed(-121,32);
				when 2993 => sin_data_int <= to_signed(-993,32); cos_data_int <= to_signed(-119,32);
				when 2994 => sin_data_int <= to_signed(-993,32); cos_data_int <= to_signed(-118,32);
				when 2995 => sin_data_int <= to_signed(-993,32); cos_data_int <= to_signed(-116,32);
				when 2996 => sin_data_int <= to_signed(-993,32); cos_data_int <= to_signed(-115,32);
				when 2997 => sin_data_int <= to_signed(-993,32); cos_data_int <= to_signed(-113,32);
				when 2998 => sin_data_int <= to_signed(-994,32); cos_data_int <= to_signed(-112,32);
				when 2999 => sin_data_int <= to_signed(-994,32); cos_data_int <= to_signed(-110,32);
				when 3000 => sin_data_int <= to_signed(-994,32); cos_data_int <= to_signed(-109,32);
				when 3001 => sin_data_int <= to_signed(-994,32); cos_data_int <= to_signed(-107,32);
				when 3002 => sin_data_int <= to_signed(-994,32); cos_data_int <= to_signed(-106,32);
				when 3003 => sin_data_int <= to_signed(-994,32); cos_data_int <= to_signed(-104,32);
				when 3004 => sin_data_int <= to_signed(-995,32); cos_data_int <= to_signed(-103,32);
				when 3005 => sin_data_int <= to_signed(-995,32); cos_data_int <= to_signed(-101,32);
				when 3006 => sin_data_int <= to_signed(-995,32); cos_data_int <= to_signed(-100,32);
				when 3007 => sin_data_int <= to_signed(-995,32); cos_data_int <= to_signed(-98,32);
				when 3008 => sin_data_int <= to_signed(-995,32); cos_data_int <= to_signed(-96,32);
				when 3009 => sin_data_int <= to_signed(-995,32); cos_data_int <= to_signed(-95,32);
				when 3010 => sin_data_int <= to_signed(-995,32); cos_data_int <= to_signed(-93,32);
				when 3011 => sin_data_int <= to_signed(-996,32); cos_data_int <= to_signed(-92,32);
				when 3012 => sin_data_int <= to_signed(-996,32); cos_data_int <= to_signed(-90,32);
				when 3013 => sin_data_int <= to_signed(-996,32); cos_data_int <= to_signed(-89,32);
				when 3014 => sin_data_int <= to_signed(-996,32); cos_data_int <= to_signed(-87,32);
				when 3015 => sin_data_int <= to_signed(-996,32); cos_data_int <= to_signed(-86,32);
				when 3016 => sin_data_int <= to_signed(-996,32); cos_data_int <= to_signed(-84,32);
				when 3017 => sin_data_int <= to_signed(-996,32); cos_data_int <= to_signed(-83,32);
				when 3018 => sin_data_int <= to_signed(-997,32); cos_data_int <= to_signed(-81,32);
				when 3019 => sin_data_int <= to_signed(-997,32); cos_data_int <= to_signed(-80,32);
				when 3020 => sin_data_int <= to_signed(-997,32); cos_data_int <= to_signed(-78,32);
				when 3021 => sin_data_int <= to_signed(-997,32); cos_data_int <= to_signed(-77,32);
				when 3022 => sin_data_int <= to_signed(-997,32); cos_data_int <= to_signed(-75,32);
				when 3023 => sin_data_int <= to_signed(-997,32); cos_data_int <= to_signed(-74,32);
				when 3024 => sin_data_int <= to_signed(-997,32); cos_data_int <= to_signed(-72,32);
				when 3025 => sin_data_int <= to_signed(-997,32); cos_data_int <= to_signed(-71,32);
				when 3026 => sin_data_int <= to_signed(-998,32); cos_data_int <= to_signed(-69,32);
				when 3027 => sin_data_int <= to_signed(-998,32); cos_data_int <= to_signed(-67,32);
				when 3028 => sin_data_int <= to_signed(-998,32); cos_data_int <= to_signed(-66,32);
				when 3029 => sin_data_int <= to_signed(-998,32); cos_data_int <= to_signed(-64,32);
				when 3030 => sin_data_int <= to_signed(-998,32); cos_data_int <= to_signed(-63,32);
				when 3031 => sin_data_int <= to_signed(-998,32); cos_data_int <= to_signed(-61,32);
				when 3032 => sin_data_int <= to_signed(-998,32); cos_data_int <= to_signed(-60,32);
				when 3033 => sin_data_int <= to_signed(-998,32); cos_data_int <= to_signed(-58,32);
				when 3034 => sin_data_int <= to_signed(-998,32); cos_data_int <= to_signed(-57,32);
				when 3035 => sin_data_int <= to_signed(-998,32); cos_data_int <= to_signed(-55,32);
				when 3036 => sin_data_int <= to_signed(-998,32); cos_data_int <= to_signed(-54,32);
				when 3037 => sin_data_int <= to_signed(-999,32); cos_data_int <= to_signed(-52,32);
				when 3038 => sin_data_int <= to_signed(-999,32); cos_data_int <= to_signed(-51,32);
				when 3039 => sin_data_int <= to_signed(-999,32); cos_data_int <= to_signed(-49,32);
				when 3040 => sin_data_int <= to_signed(-999,32); cos_data_int <= to_signed(-48,32);
				when 3041 => sin_data_int <= to_signed(-999,32); cos_data_int <= to_signed(-46,32);
				when 3042 => sin_data_int <= to_signed(-999,32); cos_data_int <= to_signed(-44,32);
				when 3043 => sin_data_int <= to_signed(-999,32); cos_data_int <= to_signed(-43,32);
				when 3044 => sin_data_int <= to_signed(-999,32); cos_data_int <= to_signed(-41,32);
				when 3045 => sin_data_int <= to_signed(-999,32); cos_data_int <= to_signed(-40,32);
				when 3046 => sin_data_int <= to_signed(-999,32); cos_data_int <= to_signed(-38,32);
				when 3047 => sin_data_int <= to_signed(-999,32); cos_data_int <= to_signed(-37,32);
				when 3048 => sin_data_int <= to_signed(-999,32); cos_data_int <= to_signed(-35,32);
				when 3049 => sin_data_int <= to_signed(-999,32); cos_data_int <= to_signed(-34,32);
				when 3050 => sin_data_int <= to_signed(-999,32); cos_data_int <= to_signed(-32,32);
				when 3051 => sin_data_int <= to_signed(-999,32); cos_data_int <= to_signed(-31,32);
				when 3052 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(-29,32);
				when 3053 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(-28,32);
				when 3054 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(-26,32);
				when 3055 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(-25,32);
				when 3056 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(-23,32);
				when 3057 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(-21,32);
				when 3058 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(-20,32);
				when 3059 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(-18,32);
				when 3060 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(-17,32);
				when 3061 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(-15,32);
				when 3062 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(-14,32);
				when 3063 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(-12,32);
				when 3064 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(-11,32);
				when 3065 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(-9,32);
				when 3066 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(-8,32);
				when 3067 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(-6,32);
				when 3068 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(-5,32);
				when 3069 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(-3,32);
				when 3070 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(-2,32);
				when 3071 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(0,32);
				when 3072 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(2,32);
				when 3073 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(3,32);
				when 3074 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(5,32);
				when 3075 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(6,32);
				when 3076 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(8,32);
				when 3077 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(9,32);
				when 3078 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(11,32);
				when 3079 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(12,32);
				when 3080 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(14,32);
				when 3081 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(15,32);
				when 3082 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(17,32);
				when 3083 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(18,32);
				when 3084 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(20,32);
				when 3085 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(21,32);
				when 3086 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(23,32);
				when 3087 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(25,32);
				when 3088 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(26,32);
				when 3089 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(28,32);
				when 3090 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(29,32);
				when 3091 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(31,32);
				when 3092 => sin_data_int <= to_signed(-1000,32); cos_data_int <= to_signed(32,32);
				when 3093 => sin_data_int <= to_signed(-999,32); cos_data_int <= to_signed(34,32);
				when 3094 => sin_data_int <= to_signed(-999,32); cos_data_int <= to_signed(35,32);
				when 3095 => sin_data_int <= to_signed(-999,32); cos_data_int <= to_signed(37,32);
				when 3096 => sin_data_int <= to_signed(-999,32); cos_data_int <= to_signed(38,32);
				when 3097 => sin_data_int <= to_signed(-999,32); cos_data_int <= to_signed(40,32);
				when 3098 => sin_data_int <= to_signed(-999,32); cos_data_int <= to_signed(41,32);
				when 3099 => sin_data_int <= to_signed(-999,32); cos_data_int <= to_signed(43,32);
				when 3100 => sin_data_int <= to_signed(-999,32); cos_data_int <= to_signed(44,32);
				when 3101 => sin_data_int <= to_signed(-999,32); cos_data_int <= to_signed(46,32);
				when 3102 => sin_data_int <= to_signed(-999,32); cos_data_int <= to_signed(48,32);
				when 3103 => sin_data_int <= to_signed(-999,32); cos_data_int <= to_signed(49,32);
				when 3104 => sin_data_int <= to_signed(-999,32); cos_data_int <= to_signed(51,32);
				when 3105 => sin_data_int <= to_signed(-999,32); cos_data_int <= to_signed(52,32);
				when 3106 => sin_data_int <= to_signed(-999,32); cos_data_int <= to_signed(54,32);
				when 3107 => sin_data_int <= to_signed(-999,32); cos_data_int <= to_signed(55,32);
				when 3108 => sin_data_int <= to_signed(-998,32); cos_data_int <= to_signed(57,32);
				when 3109 => sin_data_int <= to_signed(-998,32); cos_data_int <= to_signed(58,32);
				when 3110 => sin_data_int <= to_signed(-998,32); cos_data_int <= to_signed(60,32);
				when 3111 => sin_data_int <= to_signed(-998,32); cos_data_int <= to_signed(61,32);
				when 3112 => sin_data_int <= to_signed(-998,32); cos_data_int <= to_signed(63,32);
				when 3113 => sin_data_int <= to_signed(-998,32); cos_data_int <= to_signed(64,32);
				when 3114 => sin_data_int <= to_signed(-998,32); cos_data_int <= to_signed(66,32);
				when 3115 => sin_data_int <= to_signed(-998,32); cos_data_int <= to_signed(67,32);
				when 3116 => sin_data_int <= to_signed(-998,32); cos_data_int <= to_signed(69,32);
				when 3117 => sin_data_int <= to_signed(-998,32); cos_data_int <= to_signed(71,32);
				when 3118 => sin_data_int <= to_signed(-998,32); cos_data_int <= to_signed(72,32);
				when 3119 => sin_data_int <= to_signed(-997,32); cos_data_int <= to_signed(74,32);
				when 3120 => sin_data_int <= to_signed(-997,32); cos_data_int <= to_signed(75,32);
				when 3121 => sin_data_int <= to_signed(-997,32); cos_data_int <= to_signed(77,32);
				when 3122 => sin_data_int <= to_signed(-997,32); cos_data_int <= to_signed(78,32);
				when 3123 => sin_data_int <= to_signed(-997,32); cos_data_int <= to_signed(80,32);
				when 3124 => sin_data_int <= to_signed(-997,32); cos_data_int <= to_signed(81,32);
				when 3125 => sin_data_int <= to_signed(-997,32); cos_data_int <= to_signed(83,32);
				when 3126 => sin_data_int <= to_signed(-997,32); cos_data_int <= to_signed(84,32);
				when 3127 => sin_data_int <= to_signed(-996,32); cos_data_int <= to_signed(86,32);
				when 3128 => sin_data_int <= to_signed(-996,32); cos_data_int <= to_signed(87,32);
				when 3129 => sin_data_int <= to_signed(-996,32); cos_data_int <= to_signed(89,32);
				when 3130 => sin_data_int <= to_signed(-996,32); cos_data_int <= to_signed(90,32);
				when 3131 => sin_data_int <= to_signed(-996,32); cos_data_int <= to_signed(92,32);
				when 3132 => sin_data_int <= to_signed(-996,32); cos_data_int <= to_signed(93,32);
				when 3133 => sin_data_int <= to_signed(-996,32); cos_data_int <= to_signed(95,32);
				when 3134 => sin_data_int <= to_signed(-995,32); cos_data_int <= to_signed(96,32);
				when 3135 => sin_data_int <= to_signed(-995,32); cos_data_int <= to_signed(98,32);
				when 3136 => sin_data_int <= to_signed(-995,32); cos_data_int <= to_signed(100,32);
				when 3137 => sin_data_int <= to_signed(-995,32); cos_data_int <= to_signed(101,32);
				when 3138 => sin_data_int <= to_signed(-995,32); cos_data_int <= to_signed(103,32);
				when 3139 => sin_data_int <= to_signed(-995,32); cos_data_int <= to_signed(104,32);
				when 3140 => sin_data_int <= to_signed(-995,32); cos_data_int <= to_signed(106,32);
				when 3141 => sin_data_int <= to_signed(-994,32); cos_data_int <= to_signed(107,32);
				when 3142 => sin_data_int <= to_signed(-994,32); cos_data_int <= to_signed(109,32);
				when 3143 => sin_data_int <= to_signed(-994,32); cos_data_int <= to_signed(110,32);
				when 3144 => sin_data_int <= to_signed(-994,32); cos_data_int <= to_signed(112,32);
				when 3145 => sin_data_int <= to_signed(-994,32); cos_data_int <= to_signed(113,32);
				when 3146 => sin_data_int <= to_signed(-994,32); cos_data_int <= to_signed(115,32);
				when 3147 => sin_data_int <= to_signed(-993,32); cos_data_int <= to_signed(116,32);
				when 3148 => sin_data_int <= to_signed(-993,32); cos_data_int <= to_signed(118,32);
				when 3149 => sin_data_int <= to_signed(-993,32); cos_data_int <= to_signed(119,32);
				when 3150 => sin_data_int <= to_signed(-993,32); cos_data_int <= to_signed(121,32);
				when 3151 => sin_data_int <= to_signed(-993,32); cos_data_int <= to_signed(122,32);
				when 3152 => sin_data_int <= to_signed(-992,32); cos_data_int <= to_signed(124,32);
				when 3153 => sin_data_int <= to_signed(-992,32); cos_data_int <= to_signed(125,32);
				when 3154 => sin_data_int <= to_signed(-992,32); cos_data_int <= to_signed(127,32);
				when 3155 => sin_data_int <= to_signed(-992,32); cos_data_int <= to_signed(128,32);
				when 3156 => sin_data_int <= to_signed(-992,32); cos_data_int <= to_signed(130,32);
				when 3157 => sin_data_int <= to_signed(-992,32); cos_data_int <= to_signed(132,32);
				when 3158 => sin_data_int <= to_signed(-991,32); cos_data_int <= to_signed(133,32);
				when 3159 => sin_data_int <= to_signed(-991,32); cos_data_int <= to_signed(135,32);
				when 3160 => sin_data_int <= to_signed(-991,32); cos_data_int <= to_signed(136,32);
				when 3161 => sin_data_int <= to_signed(-991,32); cos_data_int <= to_signed(138,32);
				when 3162 => sin_data_int <= to_signed(-990,32); cos_data_int <= to_signed(139,32);
				when 3163 => sin_data_int <= to_signed(-990,32); cos_data_int <= to_signed(141,32);
				when 3164 => sin_data_int <= to_signed(-990,32); cos_data_int <= to_signed(142,32);
				when 3165 => sin_data_int <= to_signed(-990,32); cos_data_int <= to_signed(144,32);
				when 3166 => sin_data_int <= to_signed(-990,32); cos_data_int <= to_signed(145,32);
				when 3167 => sin_data_int <= to_signed(-989,32); cos_data_int <= to_signed(147,32);
				when 3168 => sin_data_int <= to_signed(-989,32); cos_data_int <= to_signed(148,32);
				when 3169 => sin_data_int <= to_signed(-989,32); cos_data_int <= to_signed(150,32);
				when 3170 => sin_data_int <= to_signed(-989,32); cos_data_int <= to_signed(151,32);
				when 3171 => sin_data_int <= to_signed(-988,32); cos_data_int <= to_signed(153,32);
				when 3172 => sin_data_int <= to_signed(-988,32); cos_data_int <= to_signed(154,32);
				when 3173 => sin_data_int <= to_signed(-988,32); cos_data_int <= to_signed(156,32);
				when 3174 => sin_data_int <= to_signed(-988,32); cos_data_int <= to_signed(157,32);
				when 3175 => sin_data_int <= to_signed(-988,32); cos_data_int <= to_signed(159,32);
				when 3176 => sin_data_int <= to_signed(-987,32); cos_data_int <= to_signed(160,32);
				when 3177 => sin_data_int <= to_signed(-987,32); cos_data_int <= to_signed(162,32);
				when 3178 => sin_data_int <= to_signed(-987,32); cos_data_int <= to_signed(163,32);
				when 3179 => sin_data_int <= to_signed(-987,32); cos_data_int <= to_signed(165,32);
				when 3180 => sin_data_int <= to_signed(-986,32); cos_data_int <= to_signed(166,32);
				when 3181 => sin_data_int <= to_signed(-986,32); cos_data_int <= to_signed(168,32);
				when 3182 => sin_data_int <= to_signed(-986,32); cos_data_int <= to_signed(169,32);
				when 3183 => sin_data_int <= to_signed(-986,32); cos_data_int <= to_signed(171,32);
				when 3184 => sin_data_int <= to_signed(-985,32); cos_data_int <= to_signed(172,32);
				when 3185 => sin_data_int <= to_signed(-985,32); cos_data_int <= to_signed(174,32);
				when 3186 => sin_data_int <= to_signed(-985,32); cos_data_int <= to_signed(175,32);
				when 3187 => sin_data_int <= to_signed(-984,32); cos_data_int <= to_signed(177,32);
				when 3188 => sin_data_int <= to_signed(-984,32); cos_data_int <= to_signed(179,32);
				when 3189 => sin_data_int <= to_signed(-984,32); cos_data_int <= to_signed(180,32);
				when 3190 => sin_data_int <= to_signed(-984,32); cos_data_int <= to_signed(182,32);
				when 3191 => sin_data_int <= to_signed(-983,32); cos_data_int <= to_signed(183,32);
				when 3192 => sin_data_int <= to_signed(-983,32); cos_data_int <= to_signed(185,32);
				when 3193 => sin_data_int <= to_signed(-983,32); cos_data_int <= to_signed(186,32);
				when 3194 => sin_data_int <= to_signed(-983,32); cos_data_int <= to_signed(188,32);
				when 3195 => sin_data_int <= to_signed(-982,32); cos_data_int <= to_signed(189,32);
				when 3196 => sin_data_int <= to_signed(-982,32); cos_data_int <= to_signed(191,32);
				when 3197 => sin_data_int <= to_signed(-982,32); cos_data_int <= to_signed(192,32);
				when 3198 => sin_data_int <= to_signed(-981,32); cos_data_int <= to_signed(194,32);
				when 3199 => sin_data_int <= to_signed(-981,32); cos_data_int <= to_signed(195,32);
				when 3200 => sin_data_int <= to_signed(-981,32); cos_data_int <= to_signed(197,32);
				when 3201 => sin_data_int <= to_signed(-980,32); cos_data_int <= to_signed(198,32);
				when 3202 => sin_data_int <= to_signed(-980,32); cos_data_int <= to_signed(200,32);
				when 3203 => sin_data_int <= to_signed(-980,32); cos_data_int <= to_signed(201,32);
				when 3204 => sin_data_int <= to_signed(-980,32); cos_data_int <= to_signed(203,32);
				when 3205 => sin_data_int <= to_signed(-979,32); cos_data_int <= to_signed(204,32);
				when 3206 => sin_data_int <= to_signed(-979,32); cos_data_int <= to_signed(206,32);
				when 3207 => sin_data_int <= to_signed(-979,32); cos_data_int <= to_signed(207,32);
				when 3208 => sin_data_int <= to_signed(-978,32); cos_data_int <= to_signed(209,32);
				when 3209 => sin_data_int <= to_signed(-978,32); cos_data_int <= to_signed(210,32);
				when 3210 => sin_data_int <= to_signed(-978,32); cos_data_int <= to_signed(212,32);
				when 3211 => sin_data_int <= to_signed(-977,32); cos_data_int <= to_signed(213,32);
				when 3212 => sin_data_int <= to_signed(-977,32); cos_data_int <= to_signed(215,32);
				when 3213 => sin_data_int <= to_signed(-977,32); cos_data_int <= to_signed(216,32);
				when 3214 => sin_data_int <= to_signed(-976,32); cos_data_int <= to_signed(218,32);
				when 3215 => sin_data_int <= to_signed(-976,32); cos_data_int <= to_signed(219,32);
				when 3216 => sin_data_int <= to_signed(-976,32); cos_data_int <= to_signed(221,32);
				when 3217 => sin_data_int <= to_signed(-975,32); cos_data_int <= to_signed(222,32);
				when 3218 => sin_data_int <= to_signed(-975,32); cos_data_int <= to_signed(224,32);
				when 3219 => sin_data_int <= to_signed(-975,32); cos_data_int <= to_signed(225,32);
				when 3220 => sin_data_int <= to_signed(-974,32); cos_data_int <= to_signed(227,32);
				when 3221 => sin_data_int <= to_signed(-974,32); cos_data_int <= to_signed(228,32);
				when 3222 => sin_data_int <= to_signed(-974,32); cos_data_int <= to_signed(230,32);
				when 3223 => sin_data_int <= to_signed(-973,32); cos_data_int <= to_signed(231,32);
				when 3224 => sin_data_int <= to_signed(-973,32); cos_data_int <= to_signed(233,32);
				when 3225 => sin_data_int <= to_signed(-973,32); cos_data_int <= to_signed(234,32);
				when 3226 => sin_data_int <= to_signed(-972,32); cos_data_int <= to_signed(236,32);
				when 3227 => sin_data_int <= to_signed(-972,32); cos_data_int <= to_signed(237,32);
				when 3228 => sin_data_int <= to_signed(-972,32); cos_data_int <= to_signed(239,32);
				when 3229 => sin_data_int <= to_signed(-971,32); cos_data_int <= to_signed(240,32);
				when 3230 => sin_data_int <= to_signed(-971,32); cos_data_int <= to_signed(241,32);
				when 3231 => sin_data_int <= to_signed(-970,32); cos_data_int <= to_signed(243,32);
				when 3232 => sin_data_int <= to_signed(-970,32); cos_data_int <= to_signed(244,32);
				when 3233 => sin_data_int <= to_signed(-970,32); cos_data_int <= to_signed(246,32);
				when 3234 => sin_data_int <= to_signed(-969,32); cos_data_int <= to_signed(247,32);
				when 3235 => sin_data_int <= to_signed(-969,32); cos_data_int <= to_signed(249,32);
				when 3236 => sin_data_int <= to_signed(-969,32); cos_data_int <= to_signed(250,32);
				when 3237 => sin_data_int <= to_signed(-968,32); cos_data_int <= to_signed(252,32);
				when 3238 => sin_data_int <= to_signed(-968,32); cos_data_int <= to_signed(253,32);
				when 3239 => sin_data_int <= to_signed(-967,32); cos_data_int <= to_signed(255,32);
				when 3240 => sin_data_int <= to_signed(-967,32); cos_data_int <= to_signed(256,32);
				when 3241 => sin_data_int <= to_signed(-967,32); cos_data_int <= to_signed(258,32);
				when 3242 => sin_data_int <= to_signed(-966,32); cos_data_int <= to_signed(259,32);
				when 3243 => sin_data_int <= to_signed(-966,32); cos_data_int <= to_signed(261,32);
				when 3244 => sin_data_int <= to_signed(-965,32); cos_data_int <= to_signed(262,32);
				when 3245 => sin_data_int <= to_signed(-965,32); cos_data_int <= to_signed(264,32);
				when 3246 => sin_data_int <= to_signed(-965,32); cos_data_int <= to_signed(265,32);
				when 3247 => sin_data_int <= to_signed(-964,32); cos_data_int <= to_signed(267,32);
				when 3248 => sin_data_int <= to_signed(-964,32); cos_data_int <= to_signed(268,32);
				when 3249 => sin_data_int <= to_signed(-963,32); cos_data_int <= to_signed(270,32);
				when 3250 => sin_data_int <= to_signed(-963,32); cos_data_int <= to_signed(271,32);
				when 3251 => sin_data_int <= to_signed(-963,32); cos_data_int <= to_signed(273,32);
				when 3252 => sin_data_int <= to_signed(-962,32); cos_data_int <= to_signed(274,32);
				when 3253 => sin_data_int <= to_signed(-962,32); cos_data_int <= to_signed(276,32);
				when 3254 => sin_data_int <= to_signed(-961,32); cos_data_int <= to_signed(277,32);
				when 3255 => sin_data_int <= to_signed(-961,32); cos_data_int <= to_signed(279,32);
				when 3256 => sin_data_int <= to_signed(-960,32); cos_data_int <= to_signed(280,32);
				when 3257 => sin_data_int <= to_signed(-960,32); cos_data_int <= to_signed(281,32);
				when 3258 => sin_data_int <= to_signed(-960,32); cos_data_int <= to_signed(283,32);
				when 3259 => sin_data_int <= to_signed(-959,32); cos_data_int <= to_signed(284,32);
				when 3260 => sin_data_int <= to_signed(-959,32); cos_data_int <= to_signed(286,32);
				when 3261 => sin_data_int <= to_signed(-958,32); cos_data_int <= to_signed(287,32);
				when 3262 => sin_data_int <= to_signed(-958,32); cos_data_int <= to_signed(289,32);
				when 3263 => sin_data_int <= to_signed(-957,32); cos_data_int <= to_signed(290,32);
				when 3264 => sin_data_int <= to_signed(-957,32); cos_data_int <= to_signed(292,32);
				when 3265 => sin_data_int <= to_signed(-956,32); cos_data_int <= to_signed(293,32);
				when 3266 => sin_data_int <= to_signed(-956,32); cos_data_int <= to_signed(295,32);
				when 3267 => sin_data_int <= to_signed(-956,32); cos_data_int <= to_signed(296,32);
				when 3268 => sin_data_int <= to_signed(-955,32); cos_data_int <= to_signed(298,32);
				when 3269 => sin_data_int <= to_signed(-955,32); cos_data_int <= to_signed(299,32);
				when 3270 => sin_data_int <= to_signed(-954,32); cos_data_int <= to_signed(301,32);
				when 3271 => sin_data_int <= to_signed(-954,32); cos_data_int <= to_signed(302,32);
				when 3272 => sin_data_int <= to_signed(-953,32); cos_data_int <= to_signed(303,32);
				when 3273 => sin_data_int <= to_signed(-953,32); cos_data_int <= to_signed(305,32);
				when 3274 => sin_data_int <= to_signed(-952,32); cos_data_int <= to_signed(306,32);
				when 3275 => sin_data_int <= to_signed(-952,32); cos_data_int <= to_signed(308,32);
				when 3276 => sin_data_int <= to_signed(-951,32); cos_data_int <= to_signed(309,32);
				when 3277 => sin_data_int <= to_signed(-951,32); cos_data_int <= to_signed(311,32);
				when 3278 => sin_data_int <= to_signed(-950,32); cos_data_int <= to_signed(312,32);
				when 3279 => sin_data_int <= to_signed(-950,32); cos_data_int <= to_signed(314,32);
				when 3280 => sin_data_int <= to_signed(-950,32); cos_data_int <= to_signed(315,32);
				when 3281 => sin_data_int <= to_signed(-949,32); cos_data_int <= to_signed(317,32);
				when 3282 => sin_data_int <= to_signed(-949,32); cos_data_int <= to_signed(318,32);
				when 3283 => sin_data_int <= to_signed(-948,32); cos_data_int <= to_signed(320,32);
				when 3284 => sin_data_int <= to_signed(-948,32); cos_data_int <= to_signed(321,32);
				when 3285 => sin_data_int <= to_signed(-947,32); cos_data_int <= to_signed(322,32);
				when 3286 => sin_data_int <= to_signed(-947,32); cos_data_int <= to_signed(324,32);
				when 3287 => sin_data_int <= to_signed(-946,32); cos_data_int <= to_signed(325,32);
				when 3288 => sin_data_int <= to_signed(-946,32); cos_data_int <= to_signed(327,32);
				when 3289 => sin_data_int <= to_signed(-945,32); cos_data_int <= to_signed(328,32);
				when 3290 => sin_data_int <= to_signed(-945,32); cos_data_int <= to_signed(330,32);
				when 3291 => sin_data_int <= to_signed(-944,32); cos_data_int <= to_signed(331,32);
				when 3292 => sin_data_int <= to_signed(-944,32); cos_data_int <= to_signed(333,32);
				when 3293 => sin_data_int <= to_signed(-943,32); cos_data_int <= to_signed(334,32);
				when 3294 => sin_data_int <= to_signed(-943,32); cos_data_int <= to_signed(335,32);
				when 3295 => sin_data_int <= to_signed(-942,32); cos_data_int <= to_signed(337,32);
				when 3296 => sin_data_int <= to_signed(-942,32); cos_data_int <= to_signed(338,32);
				when 3297 => sin_data_int <= to_signed(-941,32); cos_data_int <= to_signed(340,32);
				when 3298 => sin_data_int <= to_signed(-941,32); cos_data_int <= to_signed(341,32);
				when 3299 => sin_data_int <= to_signed(-940,32); cos_data_int <= to_signed(343,32);
				when 3300 => sin_data_int <= to_signed(-939,32); cos_data_int <= to_signed(344,32);
				when 3301 => sin_data_int <= to_signed(-939,32); cos_data_int <= to_signed(346,32);
				when 3302 => sin_data_int <= to_signed(-938,32); cos_data_int <= to_signed(347,32);
				when 3303 => sin_data_int <= to_signed(-938,32); cos_data_int <= to_signed(348,32);
				when 3304 => sin_data_int <= to_signed(-937,32); cos_data_int <= to_signed(350,32);
				when 3305 => sin_data_int <= to_signed(-937,32); cos_data_int <= to_signed(351,32);
				when 3306 => sin_data_int <= to_signed(-936,32); cos_data_int <= to_signed(353,32);
				when 3307 => sin_data_int <= to_signed(-936,32); cos_data_int <= to_signed(354,32);
				when 3308 => sin_data_int <= to_signed(-935,32); cos_data_int <= to_signed(356,32);
				when 3309 => sin_data_int <= to_signed(-935,32); cos_data_int <= to_signed(357,32);
				when 3310 => sin_data_int <= to_signed(-934,32); cos_data_int <= to_signed(358,32);
				when 3311 => sin_data_int <= to_signed(-934,32); cos_data_int <= to_signed(360,32);
				when 3312 => sin_data_int <= to_signed(-933,32); cos_data_int <= to_signed(361,32);
				when 3313 => sin_data_int <= to_signed(-932,32); cos_data_int <= to_signed(363,32);
				when 3314 => sin_data_int <= to_signed(-932,32); cos_data_int <= to_signed(364,32);
				when 3315 => sin_data_int <= to_signed(-931,32); cos_data_int <= to_signed(366,32);
				when 3316 => sin_data_int <= to_signed(-931,32); cos_data_int <= to_signed(367,32);
				when 3317 => sin_data_int <= to_signed(-930,32); cos_data_int <= to_signed(368,32);
				when 3318 => sin_data_int <= to_signed(-930,32); cos_data_int <= to_signed(370,32);
				when 3319 => sin_data_int <= to_signed(-929,32); cos_data_int <= to_signed(371,32);
				when 3320 => sin_data_int <= to_signed(-929,32); cos_data_int <= to_signed(373,32);
				when 3321 => sin_data_int <= to_signed(-928,32); cos_data_int <= to_signed(374,32);
				when 3322 => sin_data_int <= to_signed(-927,32); cos_data_int <= to_signed(376,32);
				when 3323 => sin_data_int <= to_signed(-927,32); cos_data_int <= to_signed(377,32);
				when 3324 => sin_data_int <= to_signed(-926,32); cos_data_int <= to_signed(378,32);
				when 3325 => sin_data_int <= to_signed(-926,32); cos_data_int <= to_signed(380,32);
				when 3326 => sin_data_int <= to_signed(-925,32); cos_data_int <= to_signed(381,32);
				when 3327 => sin_data_int <= to_signed(-924,32); cos_data_int <= to_signed(383,32);
				when 3328 => sin_data_int <= to_signed(-924,32); cos_data_int <= to_signed(384,32);
				when 3329 => sin_data_int <= to_signed(-923,32); cos_data_int <= to_signed(386,32);
				when 3330 => sin_data_int <= to_signed(-923,32); cos_data_int <= to_signed(387,32);
				when 3331 => sin_data_int <= to_signed(-922,32); cos_data_int <= to_signed(388,32);
				when 3332 => sin_data_int <= to_signed(-922,32); cos_data_int <= to_signed(390,32);
				when 3333 => sin_data_int <= to_signed(-921,32); cos_data_int <= to_signed(391,32);
				when 3334 => sin_data_int <= to_signed(-920,32); cos_data_int <= to_signed(393,32);
				when 3335 => sin_data_int <= to_signed(-920,32); cos_data_int <= to_signed(394,32);
				when 3336 => sin_data_int <= to_signed(-919,32); cos_data_int <= to_signed(395,32);
				when 3337 => sin_data_int <= to_signed(-919,32); cos_data_int <= to_signed(397,32);
				when 3338 => sin_data_int <= to_signed(-918,32); cos_data_int <= to_signed(398,32);
				when 3339 => sin_data_int <= to_signed(-917,32); cos_data_int <= to_signed(400,32);
				when 3340 => sin_data_int <= to_signed(-917,32); cos_data_int <= to_signed(401,32);
				when 3341 => sin_data_int <= to_signed(-916,32); cos_data_int <= to_signed(402,32);
				when 3342 => sin_data_int <= to_signed(-915,32); cos_data_int <= to_signed(404,32);
				when 3343 => sin_data_int <= to_signed(-915,32); cos_data_int <= to_signed(405,32);
				when 3344 => sin_data_int <= to_signed(-914,32); cos_data_int <= to_signed(407,32);
				when 3345 => sin_data_int <= to_signed(-914,32); cos_data_int <= to_signed(408,32);
				when 3346 => sin_data_int <= to_signed(-913,32); cos_data_int <= to_signed(409,32);
				when 3347 => sin_data_int <= to_signed(-912,32); cos_data_int <= to_signed(411,32);
				when 3348 => sin_data_int <= to_signed(-912,32); cos_data_int <= to_signed(412,32);
				when 3349 => sin_data_int <= to_signed(-911,32); cos_data_int <= to_signed(414,32);
				when 3350 => sin_data_int <= to_signed(-910,32); cos_data_int <= to_signed(415,32);
				when 3351 => sin_data_int <= to_signed(-910,32); cos_data_int <= to_signed(416,32);
				when 3352 => sin_data_int <= to_signed(-909,32); cos_data_int <= to_signed(418,32);
				when 3353 => sin_data_int <= to_signed(-909,32); cos_data_int <= to_signed(419,32);
				when 3354 => sin_data_int <= to_signed(-908,32); cos_data_int <= to_signed(421,32);
				when 3355 => sin_data_int <= to_signed(-907,32); cos_data_int <= to_signed(422,32);
				when 3356 => sin_data_int <= to_signed(-907,32); cos_data_int <= to_signed(423,32);
				when 3357 => sin_data_int <= to_signed(-906,32); cos_data_int <= to_signed(425,32);
				when 3358 => sin_data_int <= to_signed(-905,32); cos_data_int <= to_signed(426,32);
				when 3359 => sin_data_int <= to_signed(-905,32); cos_data_int <= to_signed(428,32);
				when 3360 => sin_data_int <= to_signed(-904,32); cos_data_int <= to_signed(429,32);
				when 3361 => sin_data_int <= to_signed(-903,32); cos_data_int <= to_signed(430,32);
				when 3362 => sin_data_int <= to_signed(-903,32); cos_data_int <= to_signed(432,32);
				when 3363 => sin_data_int <= to_signed(-902,32); cos_data_int <= to_signed(433,32);
				when 3364 => sin_data_int <= to_signed(-901,32); cos_data_int <= to_signed(434,32);
				when 3365 => sin_data_int <= to_signed(-901,32); cos_data_int <= to_signed(436,32);
				when 3366 => sin_data_int <= to_signed(-900,32); cos_data_int <= to_signed(437,32);
				when 3367 => sin_data_int <= to_signed(-899,32); cos_data_int <= to_signed(439,32);
				when 3368 => sin_data_int <= to_signed(-899,32); cos_data_int <= to_signed(440,32);
				when 3369 => sin_data_int <= to_signed(-898,32); cos_data_int <= to_signed(441,32);
				when 3370 => sin_data_int <= to_signed(-897,32); cos_data_int <= to_signed(443,32);
				when 3371 => sin_data_int <= to_signed(-897,32); cos_data_int <= to_signed(444,32);
				when 3372 => sin_data_int <= to_signed(-896,32); cos_data_int <= to_signed(445,32);
				when 3373 => sin_data_int <= to_signed(-895,32); cos_data_int <= to_signed(447,32);
				when 3374 => sin_data_int <= to_signed(-895,32); cos_data_int <= to_signed(448,32);
				when 3375 => sin_data_int <= to_signed(-894,32); cos_data_int <= to_signed(450,32);
				when 3376 => sin_data_int <= to_signed(-893,32); cos_data_int <= to_signed(451,32);
				when 3377 => sin_data_int <= to_signed(-893,32); cos_data_int <= to_signed(452,32);
				when 3378 => sin_data_int <= to_signed(-892,32); cos_data_int <= to_signed(454,32);
				when 3379 => sin_data_int <= to_signed(-891,32); cos_data_int <= to_signed(455,32);
				when 3380 => sin_data_int <= to_signed(-890,32); cos_data_int <= to_signed(456,32);
				when 3381 => sin_data_int <= to_signed(-890,32); cos_data_int <= to_signed(458,32);
				when 3382 => sin_data_int <= to_signed(-889,32); cos_data_int <= to_signed(459,32);
				when 3383 => sin_data_int <= to_signed(-888,32); cos_data_int <= to_signed(461,32);
				when 3384 => sin_data_int <= to_signed(-888,32); cos_data_int <= to_signed(462,32);
				when 3385 => sin_data_int <= to_signed(-887,32); cos_data_int <= to_signed(463,32);
				when 3386 => sin_data_int <= to_signed(-886,32); cos_data_int <= to_signed(465,32);
				when 3387 => sin_data_int <= to_signed(-886,32); cos_data_int <= to_signed(466,32);
				when 3388 => sin_data_int <= to_signed(-885,32); cos_data_int <= to_signed(467,32);
				when 3389 => sin_data_int <= to_signed(-884,32); cos_data_int <= to_signed(469,32);
				when 3390 => sin_data_int <= to_signed(-883,32); cos_data_int <= to_signed(470,32);
				when 3391 => sin_data_int <= to_signed(-883,32); cos_data_int <= to_signed(471,32);
				when 3392 => sin_data_int <= to_signed(-882,32); cos_data_int <= to_signed(473,32);
				when 3393 => sin_data_int <= to_signed(-881,32); cos_data_int <= to_signed(474,32);
				when 3394 => sin_data_int <= to_signed(-880,32); cos_data_int <= to_signed(475,32);
				when 3395 => sin_data_int <= to_signed(-880,32); cos_data_int <= to_signed(477,32);
				when 3396 => sin_data_int <= to_signed(-879,32); cos_data_int <= to_signed(478,32);
				when 3397 => sin_data_int <= to_signed(-878,32); cos_data_int <= to_signed(479,32);
				when 3398 => sin_data_int <= to_signed(-878,32); cos_data_int <= to_signed(481,32);
				when 3399 => sin_data_int <= to_signed(-877,32); cos_data_int <= to_signed(482,32);
				when 3400 => sin_data_int <= to_signed(-876,32); cos_data_int <= to_signed(484,32);
				when 3401 => sin_data_int <= to_signed(-875,32); cos_data_int <= to_signed(485,32);
				when 3402 => sin_data_int <= to_signed(-875,32); cos_data_int <= to_signed(486,32);
				when 3403 => sin_data_int <= to_signed(-874,32); cos_data_int <= to_signed(488,32);
				when 3404 => sin_data_int <= to_signed(-873,32); cos_data_int <= to_signed(489,32);
				when 3405 => sin_data_int <= to_signed(-872,32); cos_data_int <= to_signed(490,32);
				when 3406 => sin_data_int <= to_signed(-872,32); cos_data_int <= to_signed(492,32);
				when 3407 => sin_data_int <= to_signed(-871,32); cos_data_int <= to_signed(493,32);
				when 3408 => sin_data_int <= to_signed(-870,32); cos_data_int <= to_signed(494,32);
				when 3409 => sin_data_int <= to_signed(-869,32); cos_data_int <= to_signed(496,32);
				when 3410 => sin_data_int <= to_signed(-869,32); cos_data_int <= to_signed(497,32);
				when 3411 => sin_data_int <= to_signed(-868,32); cos_data_int <= to_signed(498,32);
				when 3412 => sin_data_int <= to_signed(-867,32); cos_data_int <= to_signed(500,32);
				when 3413 => sin_data_int <= to_signed(-866,32); cos_data_int <= to_signed(501,32);
				when 3414 => sin_data_int <= to_signed(-866,32); cos_data_int <= to_signed(502,32);
				when 3415 => sin_data_int <= to_signed(-865,32); cos_data_int <= to_signed(504,32);
				when 3416 => sin_data_int <= to_signed(-864,32); cos_data_int <= to_signed(505,32);
				when 3417 => sin_data_int <= to_signed(-863,32); cos_data_int <= to_signed(506,32);
				when 3418 => sin_data_int <= to_signed(-862,32); cos_data_int <= to_signed(508,32);
				when 3419 => sin_data_int <= to_signed(-862,32); cos_data_int <= to_signed(509,32);
				when 3420 => sin_data_int <= to_signed(-861,32); cos_data_int <= to_signed(510,32);
				when 3421 => sin_data_int <= to_signed(-860,32); cos_data_int <= to_signed(511,32);
				when 3422 => sin_data_int <= to_signed(-859,32); cos_data_int <= to_signed(513,32);
				when 3423 => sin_data_int <= to_signed(-859,32); cos_data_int <= to_signed(514,32);
				when 3424 => sin_data_int <= to_signed(-858,32); cos_data_int <= to_signed(515,32);
				when 3425 => sin_data_int <= to_signed(-857,32); cos_data_int <= to_signed(517,32);
				when 3426 => sin_data_int <= to_signed(-856,32); cos_data_int <= to_signed(518,32);
				when 3427 => sin_data_int <= to_signed(-855,32); cos_data_int <= to_signed(519,32);
				when 3428 => sin_data_int <= to_signed(-855,32); cos_data_int <= to_signed(521,32);
				when 3429 => sin_data_int <= to_signed(-854,32); cos_data_int <= to_signed(522,32);
				when 3430 => sin_data_int <= to_signed(-853,32); cos_data_int <= to_signed(523,32);
				when 3431 => sin_data_int <= to_signed(-852,32); cos_data_int <= to_signed(525,32);
				when 3432 => sin_data_int <= to_signed(-851,32); cos_data_int <= to_signed(526,32);
				when 3433 => sin_data_int <= to_signed(-851,32); cos_data_int <= to_signed(527,32);
				when 3434 => sin_data_int <= to_signed(-850,32); cos_data_int <= to_signed(529,32);
				when 3435 => sin_data_int <= to_signed(-849,32); cos_data_int <= to_signed(530,32);
				when 3436 => sin_data_int <= to_signed(-848,32); cos_data_int <= to_signed(531,32);
				when 3437 => sin_data_int <= to_signed(-847,32); cos_data_int <= to_signed(532,32);
				when 3438 => sin_data_int <= to_signed(-846,32); cos_data_int <= to_signed(534,32);
				when 3439 => sin_data_int <= to_signed(-846,32); cos_data_int <= to_signed(535,32);
				when 3440 => sin_data_int <= to_signed(-845,32); cos_data_int <= to_signed(536,32);
				when 3441 => sin_data_int <= to_signed(-844,32); cos_data_int <= to_signed(538,32);
				when 3442 => sin_data_int <= to_signed(-843,32); cos_data_int <= to_signed(539,32);
				when 3443 => sin_data_int <= to_signed(-842,32); cos_data_int <= to_signed(540,32);
				when 3444 => sin_data_int <= to_signed(-842,32); cos_data_int <= to_signed(541,32);
				when 3445 => sin_data_int <= to_signed(-841,32); cos_data_int <= to_signed(543,32);
				when 3446 => sin_data_int <= to_signed(-840,32); cos_data_int <= to_signed(544,32);
				when 3447 => sin_data_int <= to_signed(-839,32); cos_data_int <= to_signed(545,32);
				when 3448 => sin_data_int <= to_signed(-838,32); cos_data_int <= to_signed(547,32);
				when 3449 => sin_data_int <= to_signed(-837,32); cos_data_int <= to_signed(548,32);
				when 3450 => sin_data_int <= to_signed(-837,32); cos_data_int <= to_signed(549,32);
				when 3451 => sin_data_int <= to_signed(-836,32); cos_data_int <= to_signed(550,32);
				when 3452 => sin_data_int <= to_signed(-835,32); cos_data_int <= to_signed(552,32);
				when 3453 => sin_data_int <= to_signed(-834,32); cos_data_int <= to_signed(553,32);
				when 3454 => sin_data_int <= to_signed(-833,32); cos_data_int <= to_signed(554,32);
				when 3455 => sin_data_int <= to_signed(-832,32); cos_data_int <= to_signed(556,32);
				when 3456 => sin_data_int <= to_signed(-831,32); cos_data_int <= to_signed(557,32);
				when 3457 => sin_data_int <= to_signed(-831,32); cos_data_int <= to_signed(558,32);
				when 3458 => sin_data_int <= to_signed(-830,32); cos_data_int <= to_signed(559,32);
				when 3459 => sin_data_int <= to_signed(-829,32); cos_data_int <= to_signed(561,32);
				when 3460 => sin_data_int <= to_signed(-828,32); cos_data_int <= to_signed(562,32);
				when 3461 => sin_data_int <= to_signed(-827,32); cos_data_int <= to_signed(563,32);
				when 3462 => sin_data_int <= to_signed(-826,32); cos_data_int <= to_signed(564,32);
				when 3463 => sin_data_int <= to_signed(-825,32); cos_data_int <= to_signed(566,32);
				when 3464 => sin_data_int <= to_signed(-825,32); cos_data_int <= to_signed(567,32);
				when 3465 => sin_data_int <= to_signed(-824,32); cos_data_int <= to_signed(568,32);
				when 3466 => sin_data_int <= to_signed(-823,32); cos_data_int <= to_signed(570,32);
				when 3467 => sin_data_int <= to_signed(-822,32); cos_data_int <= to_signed(571,32);
				when 3468 => sin_data_int <= to_signed(-821,32); cos_data_int <= to_signed(572,32);
				when 3469 => sin_data_int <= to_signed(-820,32); cos_data_int <= to_signed(573,32);
				when 3470 => sin_data_int <= to_signed(-819,32); cos_data_int <= to_signed(575,32);
				when 3471 => sin_data_int <= to_signed(-818,32); cos_data_int <= to_signed(576,32);
				when 3472 => sin_data_int <= to_signed(-818,32); cos_data_int <= to_signed(577,32);
				when 3473 => sin_data_int <= to_signed(-817,32); cos_data_int <= to_signed(578,32);
				when 3474 => sin_data_int <= to_signed(-816,32); cos_data_int <= to_signed(580,32);
				when 3475 => sin_data_int <= to_signed(-815,32); cos_data_int <= to_signed(581,32);
				when 3476 => sin_data_int <= to_signed(-814,32); cos_data_int <= to_signed(582,32);
				when 3477 => sin_data_int <= to_signed(-813,32); cos_data_int <= to_signed(583,32);
				when 3478 => sin_data_int <= to_signed(-812,32); cos_data_int <= to_signed(585,32);
				when 3479 => sin_data_int <= to_signed(-811,32); cos_data_int <= to_signed(586,32);
				when 3480 => sin_data_int <= to_signed(-810,32); cos_data_int <= to_signed(587,32);
				when 3481 => sin_data_int <= to_signed(-810,32); cos_data_int <= to_signed(588,32);
				when 3482 => sin_data_int <= to_signed(-809,32); cos_data_int <= to_signed(590,32);
				when 3483 => sin_data_int <= to_signed(-808,32); cos_data_int <= to_signed(591,32);
				when 3484 => sin_data_int <= to_signed(-807,32); cos_data_int <= to_signed(592,32);
				when 3485 => sin_data_int <= to_signed(-806,32); cos_data_int <= to_signed(593,32);
				when 3486 => sin_data_int <= to_signed(-805,32); cos_data_int <= to_signed(594,32);
				when 3487 => sin_data_int <= to_signed(-804,32); cos_data_int <= to_signed(596,32);
				when 3488 => sin_data_int <= to_signed(-803,32); cos_data_int <= to_signed(597,32);
				when 3489 => sin_data_int <= to_signed(-802,32); cos_data_int <= to_signed(598,32);
				when 3490 => sin_data_int <= to_signed(-801,32); cos_data_int <= to_signed(599,32);
				when 3491 => sin_data_int <= to_signed(-800,32); cos_data_int <= to_signed(601,32);
				when 3492 => sin_data_int <= to_signed(-800,32); cos_data_int <= to_signed(602,32);
				when 3493 => sin_data_int <= to_signed(-799,32); cos_data_int <= to_signed(603,32);
				when 3494 => sin_data_int <= to_signed(-798,32); cos_data_int <= to_signed(604,32);
				when 3495 => sin_data_int <= to_signed(-797,32); cos_data_int <= to_signed(606,32);
				when 3496 => sin_data_int <= to_signed(-796,32); cos_data_int <= to_signed(607,32);
				when 3497 => sin_data_int <= to_signed(-795,32); cos_data_int <= to_signed(608,32);
				when 3498 => sin_data_int <= to_signed(-794,32); cos_data_int <= to_signed(609,32);
				when 3499 => sin_data_int <= to_signed(-793,32); cos_data_int <= to_signed(610,32);
				when 3500 => sin_data_int <= to_signed(-792,32); cos_data_int <= to_signed(612,32);
				when 3501 => sin_data_int <= to_signed(-791,32); cos_data_int <= to_signed(613,32);
				when 3502 => sin_data_int <= to_signed(-790,32); cos_data_int <= to_signed(614,32);
				when 3503 => sin_data_int <= to_signed(-789,32); cos_data_int <= to_signed(615,32);
				when 3504 => sin_data_int <= to_signed(-788,32); cos_data_int <= to_signed(616,32);
				when 3505 => sin_data_int <= to_signed(-787,32); cos_data_int <= to_signed(618,32);
				when 3506 => sin_data_int <= to_signed(-786,32); cos_data_int <= to_signed(619,32);
				when 3507 => sin_data_int <= to_signed(-786,32); cos_data_int <= to_signed(620,32);
				when 3508 => sin_data_int <= to_signed(-785,32); cos_data_int <= to_signed(621,32);
				when 3509 => sin_data_int <= to_signed(-784,32); cos_data_int <= to_signed(622,32);
				when 3510 => sin_data_int <= to_signed(-783,32); cos_data_int <= to_signed(624,32);
				when 3511 => sin_data_int <= to_signed(-782,32); cos_data_int <= to_signed(625,32);
				when 3512 => sin_data_int <= to_signed(-781,32); cos_data_int <= to_signed(626,32);
				when 3513 => sin_data_int <= to_signed(-780,32); cos_data_int <= to_signed(627,32);
				when 3514 => sin_data_int <= to_signed(-779,32); cos_data_int <= to_signed(628,32);
				when 3515 => sin_data_int <= to_signed(-778,32); cos_data_int <= to_signed(630,32);
				when 3516 => sin_data_int <= to_signed(-777,32); cos_data_int <= to_signed(631,32);
				when 3517 => sin_data_int <= to_signed(-776,32); cos_data_int <= to_signed(632,32);
				when 3518 => sin_data_int <= to_signed(-775,32); cos_data_int <= to_signed(633,32);
				when 3519 => sin_data_int <= to_signed(-774,32); cos_data_int <= to_signed(634,32);
				when 3520 => sin_data_int <= to_signed(-773,32); cos_data_int <= to_signed(636,32);
				when 3521 => sin_data_int <= to_signed(-772,32); cos_data_int <= to_signed(637,32);
				when 3522 => sin_data_int <= to_signed(-771,32); cos_data_int <= to_signed(638,32);
				when 3523 => sin_data_int <= to_signed(-770,32); cos_data_int <= to_signed(639,32);
				when 3524 => sin_data_int <= to_signed(-769,32); cos_data_int <= to_signed(640,32);
				when 3525 => sin_data_int <= to_signed(-768,32); cos_data_int <= to_signed(641,32);
				when 3526 => sin_data_int <= to_signed(-767,32); cos_data_int <= to_signed(643,32);
				when 3527 => sin_data_int <= to_signed(-766,32); cos_data_int <= to_signed(644,32);
				when 3528 => sin_data_int <= to_signed(-765,32); cos_data_int <= to_signed(645,32);
				when 3529 => sin_data_int <= to_signed(-764,32); cos_data_int <= to_signed(646,32);
				when 3530 => sin_data_int <= to_signed(-763,32); cos_data_int <= to_signed(647,32);
				when 3531 => sin_data_int <= to_signed(-762,32); cos_data_int <= to_signed(649,32);
				when 3532 => sin_data_int <= to_signed(-761,32); cos_data_int <= to_signed(650,32);
				when 3533 => sin_data_int <= to_signed(-760,32); cos_data_int <= to_signed(651,32);
				when 3534 => sin_data_int <= to_signed(-759,32); cos_data_int <= to_signed(652,32);
				when 3535 => sin_data_int <= to_signed(-758,32); cos_data_int <= to_signed(653,32);
				when 3536 => sin_data_int <= to_signed(-757,32); cos_data_int <= to_signed(654,32);
				when 3537 => sin_data_int <= to_signed(-756,32); cos_data_int <= to_signed(655,32);
				when 3538 => sin_data_int <= to_signed(-755,32); cos_data_int <= to_signed(657,32);
				when 3539 => sin_data_int <= to_signed(-754,32); cos_data_int <= to_signed(658,32);
				when 3540 => sin_data_int <= to_signed(-753,32); cos_data_int <= to_signed(659,32);
				when 3541 => sin_data_int <= to_signed(-752,32); cos_data_int <= to_signed(660,32);
				when 3542 => sin_data_int <= to_signed(-751,32); cos_data_int <= to_signed(661,32);
				when 3543 => sin_data_int <= to_signed(-750,32); cos_data_int <= to_signed(662,32);
				when 3544 => sin_data_int <= to_signed(-749,32); cos_data_int <= to_signed(664,32);
				when 3545 => sin_data_int <= to_signed(-748,32); cos_data_int <= to_signed(665,32);
				when 3546 => sin_data_int <= to_signed(-747,32); cos_data_int <= to_signed(666,32);
				when 3547 => sin_data_int <= to_signed(-746,32); cos_data_int <= to_signed(667,32);
				when 3548 => sin_data_int <= to_signed(-745,32); cos_data_int <= to_signed(668,32);
				when 3549 => sin_data_int <= to_signed(-744,32); cos_data_int <= to_signed(669,32);
				when 3550 => sin_data_int <= to_signed(-743,32); cos_data_int <= to_signed(670,32);
				when 3551 => sin_data_int <= to_signed(-742,32); cos_data_int <= to_signed(672,32);
				when 3552 => sin_data_int <= to_signed(-741,32); cos_data_int <= to_signed(673,32);
				when 3553 => sin_data_int <= to_signed(-740,32); cos_data_int <= to_signed(674,32);
				when 3554 => sin_data_int <= to_signed(-739,32); cos_data_int <= to_signed(675,32);
				when 3555 => sin_data_int <= to_signed(-738,32); cos_data_int <= to_signed(676,32);
				when 3556 => sin_data_int <= to_signed(-737,32); cos_data_int <= to_signed(677,32);
				when 3557 => sin_data_int <= to_signed(-736,32); cos_data_int <= to_signed(678,32);
				when 3558 => sin_data_int <= to_signed(-735,32); cos_data_int <= to_signed(679,32);
				when 3559 => sin_data_int <= to_signed(-734,32); cos_data_int <= to_signed(681,32);
				when 3560 => sin_data_int <= to_signed(-733,32); cos_data_int <= to_signed(682,32);
				when 3561 => sin_data_int <= to_signed(-732,32); cos_data_int <= to_signed(683,32);
				when 3562 => sin_data_int <= to_signed(-731,32); cos_data_int <= to_signed(684,32);
				when 3563 => sin_data_int <= to_signed(-730,32); cos_data_int <= to_signed(685,32);
				when 3564 => sin_data_int <= to_signed(-728,32); cos_data_int <= to_signed(686,32);
				when 3565 => sin_data_int <= to_signed(-727,32); cos_data_int <= to_signed(687,32);
				when 3566 => sin_data_int <= to_signed(-726,32); cos_data_int <= to_signed(688,32);
				when 3567 => sin_data_int <= to_signed(-725,32); cos_data_int <= to_signed(690,32);
				when 3568 => sin_data_int <= to_signed(-724,32); cos_data_int <= to_signed(691,32);
				when 3569 => sin_data_int <= to_signed(-723,32); cos_data_int <= to_signed(692,32);
				when 3570 => sin_data_int <= to_signed(-722,32); cos_data_int <= to_signed(693,32);
				when 3571 => sin_data_int <= to_signed(-721,32); cos_data_int <= to_signed(694,32);
				when 3572 => sin_data_int <= to_signed(-720,32); cos_data_int <= to_signed(695,32);
				when 3573 => sin_data_int <= to_signed(-719,32); cos_data_int <= to_signed(696,32);
				when 3574 => sin_data_int <= to_signed(-718,32); cos_data_int <= to_signed(697,32);
				when 3575 => sin_data_int <= to_signed(-717,32); cos_data_int <= to_signed(698,32);
				when 3576 => sin_data_int <= to_signed(-716,32); cos_data_int <= to_signed(699,32);
				when 3577 => sin_data_int <= to_signed(-715,32); cos_data_int <= to_signed(701,32);
				when 3578 => sin_data_int <= to_signed(-714,32); cos_data_int <= to_signed(702,32);
				when 3579 => sin_data_int <= to_signed(-713,32); cos_data_int <= to_signed(703,32);
				when 3580 => sin_data_int <= to_signed(-711,32); cos_data_int <= to_signed(704,32);
				when 3581 => sin_data_int <= to_signed(-710,32); cos_data_int <= to_signed(705,32);
				when 3582 => sin_data_int <= to_signed(-709,32); cos_data_int <= to_signed(706,32);
				when 3583 => sin_data_int <= to_signed(-708,32); cos_data_int <= to_signed(707,32);
				when 3584 => sin_data_int <= to_signed(-707,32); cos_data_int <= to_signed(708,32);
				when 3585 => sin_data_int <= to_signed(-706,32); cos_data_int <= to_signed(709,32);
				when 3586 => sin_data_int <= to_signed(-705,32); cos_data_int <= to_signed(710,32);
				when 3587 => sin_data_int <= to_signed(-704,32); cos_data_int <= to_signed(711,32);
				when 3588 => sin_data_int <= to_signed(-703,32); cos_data_int <= to_signed(713,32);
				when 3589 => sin_data_int <= to_signed(-702,32); cos_data_int <= to_signed(714,32);
				when 3590 => sin_data_int <= to_signed(-701,32); cos_data_int <= to_signed(715,32);
				when 3591 => sin_data_int <= to_signed(-699,32); cos_data_int <= to_signed(716,32);
				when 3592 => sin_data_int <= to_signed(-698,32); cos_data_int <= to_signed(717,32);
				when 3593 => sin_data_int <= to_signed(-697,32); cos_data_int <= to_signed(718,32);
				when 3594 => sin_data_int <= to_signed(-696,32); cos_data_int <= to_signed(719,32);
				when 3595 => sin_data_int <= to_signed(-695,32); cos_data_int <= to_signed(720,32);
				when 3596 => sin_data_int <= to_signed(-694,32); cos_data_int <= to_signed(721,32);
				when 3597 => sin_data_int <= to_signed(-693,32); cos_data_int <= to_signed(722,32);
				when 3598 => sin_data_int <= to_signed(-692,32); cos_data_int <= to_signed(723,32);
				when 3599 => sin_data_int <= to_signed(-691,32); cos_data_int <= to_signed(724,32);
				when 3600 => sin_data_int <= to_signed(-690,32); cos_data_int <= to_signed(725,32);
				when 3601 => sin_data_int <= to_signed(-688,32); cos_data_int <= to_signed(726,32);
				when 3602 => sin_data_int <= to_signed(-687,32); cos_data_int <= to_signed(727,32);
				when 3603 => sin_data_int <= to_signed(-686,32); cos_data_int <= to_signed(728,32);
				when 3604 => sin_data_int <= to_signed(-685,32); cos_data_int <= to_signed(730,32);
				when 3605 => sin_data_int <= to_signed(-684,32); cos_data_int <= to_signed(731,32);
				when 3606 => sin_data_int <= to_signed(-683,32); cos_data_int <= to_signed(732,32);
				when 3607 => sin_data_int <= to_signed(-682,32); cos_data_int <= to_signed(733,32);
				when 3608 => sin_data_int <= to_signed(-681,32); cos_data_int <= to_signed(734,32);
				when 3609 => sin_data_int <= to_signed(-679,32); cos_data_int <= to_signed(735,32);
				when 3610 => sin_data_int <= to_signed(-678,32); cos_data_int <= to_signed(736,32);
				when 3611 => sin_data_int <= to_signed(-677,32); cos_data_int <= to_signed(737,32);
				when 3612 => sin_data_int <= to_signed(-676,32); cos_data_int <= to_signed(738,32);
				when 3613 => sin_data_int <= to_signed(-675,32); cos_data_int <= to_signed(739,32);
				when 3614 => sin_data_int <= to_signed(-674,32); cos_data_int <= to_signed(740,32);
				when 3615 => sin_data_int <= to_signed(-673,32); cos_data_int <= to_signed(741,32);
				when 3616 => sin_data_int <= to_signed(-672,32); cos_data_int <= to_signed(742,32);
				when 3617 => sin_data_int <= to_signed(-670,32); cos_data_int <= to_signed(743,32);
				when 3618 => sin_data_int <= to_signed(-669,32); cos_data_int <= to_signed(744,32);
				when 3619 => sin_data_int <= to_signed(-668,32); cos_data_int <= to_signed(745,32);
				when 3620 => sin_data_int <= to_signed(-667,32); cos_data_int <= to_signed(746,32);
				when 3621 => sin_data_int <= to_signed(-666,32); cos_data_int <= to_signed(747,32);
				when 3622 => sin_data_int <= to_signed(-665,32); cos_data_int <= to_signed(748,32);
				when 3623 => sin_data_int <= to_signed(-664,32); cos_data_int <= to_signed(749,32);
				when 3624 => sin_data_int <= to_signed(-662,32); cos_data_int <= to_signed(750,32);
				when 3625 => sin_data_int <= to_signed(-661,32); cos_data_int <= to_signed(751,32);
				when 3626 => sin_data_int <= to_signed(-660,32); cos_data_int <= to_signed(752,32);
				when 3627 => sin_data_int <= to_signed(-659,32); cos_data_int <= to_signed(753,32);
				when 3628 => sin_data_int <= to_signed(-658,32); cos_data_int <= to_signed(754,32);
				when 3629 => sin_data_int <= to_signed(-657,32); cos_data_int <= to_signed(755,32);
				when 3630 => sin_data_int <= to_signed(-655,32); cos_data_int <= to_signed(756,32);
				when 3631 => sin_data_int <= to_signed(-654,32); cos_data_int <= to_signed(757,32);
				when 3632 => sin_data_int <= to_signed(-653,32); cos_data_int <= to_signed(758,32);
				when 3633 => sin_data_int <= to_signed(-652,32); cos_data_int <= to_signed(759,32);
				when 3634 => sin_data_int <= to_signed(-651,32); cos_data_int <= to_signed(760,32);
				when 3635 => sin_data_int <= to_signed(-650,32); cos_data_int <= to_signed(761,32);
				when 3636 => sin_data_int <= to_signed(-649,32); cos_data_int <= to_signed(762,32);
				when 3637 => sin_data_int <= to_signed(-647,32); cos_data_int <= to_signed(763,32);
				when 3638 => sin_data_int <= to_signed(-646,32); cos_data_int <= to_signed(764,32);
				when 3639 => sin_data_int <= to_signed(-645,32); cos_data_int <= to_signed(765,32);
				when 3640 => sin_data_int <= to_signed(-644,32); cos_data_int <= to_signed(766,32);
				when 3641 => sin_data_int <= to_signed(-643,32); cos_data_int <= to_signed(767,32);
				when 3642 => sin_data_int <= to_signed(-641,32); cos_data_int <= to_signed(768,32);
				when 3643 => sin_data_int <= to_signed(-640,32); cos_data_int <= to_signed(769,32);
				when 3644 => sin_data_int <= to_signed(-639,32); cos_data_int <= to_signed(770,32);
				when 3645 => sin_data_int <= to_signed(-638,32); cos_data_int <= to_signed(771,32);
				when 3646 => sin_data_int <= to_signed(-637,32); cos_data_int <= to_signed(772,32);
				when 3647 => sin_data_int <= to_signed(-636,32); cos_data_int <= to_signed(773,32);
				when 3648 => sin_data_int <= to_signed(-634,32); cos_data_int <= to_signed(774,32);
				when 3649 => sin_data_int <= to_signed(-633,32); cos_data_int <= to_signed(775,32);
				when 3650 => sin_data_int <= to_signed(-632,32); cos_data_int <= to_signed(776,32);
				when 3651 => sin_data_int <= to_signed(-631,32); cos_data_int <= to_signed(777,32);
				when 3652 => sin_data_int <= to_signed(-630,32); cos_data_int <= to_signed(778,32);
				when 3653 => sin_data_int <= to_signed(-628,32); cos_data_int <= to_signed(779,32);
				when 3654 => sin_data_int <= to_signed(-627,32); cos_data_int <= to_signed(780,32);
				when 3655 => sin_data_int <= to_signed(-626,32); cos_data_int <= to_signed(781,32);
				when 3656 => sin_data_int <= to_signed(-625,32); cos_data_int <= to_signed(782,32);
				when 3657 => sin_data_int <= to_signed(-624,32); cos_data_int <= to_signed(783,32);
				when 3658 => sin_data_int <= to_signed(-622,32); cos_data_int <= to_signed(784,32);
				when 3659 => sin_data_int <= to_signed(-621,32); cos_data_int <= to_signed(785,32);
				when 3660 => sin_data_int <= to_signed(-620,32); cos_data_int <= to_signed(786,32);
				when 3661 => sin_data_int <= to_signed(-619,32); cos_data_int <= to_signed(786,32);
				when 3662 => sin_data_int <= to_signed(-618,32); cos_data_int <= to_signed(787,32);
				when 3663 => sin_data_int <= to_signed(-616,32); cos_data_int <= to_signed(788,32);
				when 3664 => sin_data_int <= to_signed(-615,32); cos_data_int <= to_signed(789,32);
				when 3665 => sin_data_int <= to_signed(-614,32); cos_data_int <= to_signed(790,32);
				when 3666 => sin_data_int <= to_signed(-613,32); cos_data_int <= to_signed(791,32);
				when 3667 => sin_data_int <= to_signed(-612,32); cos_data_int <= to_signed(792,32);
				when 3668 => sin_data_int <= to_signed(-610,32); cos_data_int <= to_signed(793,32);
				when 3669 => sin_data_int <= to_signed(-609,32); cos_data_int <= to_signed(794,32);
				when 3670 => sin_data_int <= to_signed(-608,32); cos_data_int <= to_signed(795,32);
				when 3671 => sin_data_int <= to_signed(-607,32); cos_data_int <= to_signed(796,32);
				when 3672 => sin_data_int <= to_signed(-606,32); cos_data_int <= to_signed(797,32);
				when 3673 => sin_data_int <= to_signed(-604,32); cos_data_int <= to_signed(798,32);
				when 3674 => sin_data_int <= to_signed(-603,32); cos_data_int <= to_signed(799,32);
				when 3675 => sin_data_int <= to_signed(-602,32); cos_data_int <= to_signed(800,32);
				when 3676 => sin_data_int <= to_signed(-601,32); cos_data_int <= to_signed(800,32);
				when 3677 => sin_data_int <= to_signed(-599,32); cos_data_int <= to_signed(801,32);
				when 3678 => sin_data_int <= to_signed(-598,32); cos_data_int <= to_signed(802,32);
				when 3679 => sin_data_int <= to_signed(-597,32); cos_data_int <= to_signed(803,32);
				when 3680 => sin_data_int <= to_signed(-596,32); cos_data_int <= to_signed(804,32);
				when 3681 => sin_data_int <= to_signed(-594,32); cos_data_int <= to_signed(805,32);
				when 3682 => sin_data_int <= to_signed(-593,32); cos_data_int <= to_signed(806,32);
				when 3683 => sin_data_int <= to_signed(-592,32); cos_data_int <= to_signed(807,32);
				when 3684 => sin_data_int <= to_signed(-591,32); cos_data_int <= to_signed(808,32);
				when 3685 => sin_data_int <= to_signed(-590,32); cos_data_int <= to_signed(809,32);
				when 3686 => sin_data_int <= to_signed(-588,32); cos_data_int <= to_signed(810,32);
				when 3687 => sin_data_int <= to_signed(-587,32); cos_data_int <= to_signed(810,32);
				when 3688 => sin_data_int <= to_signed(-586,32); cos_data_int <= to_signed(811,32);
				when 3689 => sin_data_int <= to_signed(-585,32); cos_data_int <= to_signed(812,32);
				when 3690 => sin_data_int <= to_signed(-583,32); cos_data_int <= to_signed(813,32);
				when 3691 => sin_data_int <= to_signed(-582,32); cos_data_int <= to_signed(814,32);
				when 3692 => sin_data_int <= to_signed(-581,32); cos_data_int <= to_signed(815,32);
				when 3693 => sin_data_int <= to_signed(-580,32); cos_data_int <= to_signed(816,32);
				when 3694 => sin_data_int <= to_signed(-578,32); cos_data_int <= to_signed(817,32);
				when 3695 => sin_data_int <= to_signed(-577,32); cos_data_int <= to_signed(818,32);
				when 3696 => sin_data_int <= to_signed(-576,32); cos_data_int <= to_signed(818,32);
				when 3697 => sin_data_int <= to_signed(-575,32); cos_data_int <= to_signed(819,32);
				when 3698 => sin_data_int <= to_signed(-573,32); cos_data_int <= to_signed(820,32);
				when 3699 => sin_data_int <= to_signed(-572,32); cos_data_int <= to_signed(821,32);
				when 3700 => sin_data_int <= to_signed(-571,32); cos_data_int <= to_signed(822,32);
				when 3701 => sin_data_int <= to_signed(-570,32); cos_data_int <= to_signed(823,32);
				when 3702 => sin_data_int <= to_signed(-568,32); cos_data_int <= to_signed(824,32);
				when 3703 => sin_data_int <= to_signed(-567,32); cos_data_int <= to_signed(825,32);
				when 3704 => sin_data_int <= to_signed(-566,32); cos_data_int <= to_signed(825,32);
				when 3705 => sin_data_int <= to_signed(-564,32); cos_data_int <= to_signed(826,32);
				when 3706 => sin_data_int <= to_signed(-563,32); cos_data_int <= to_signed(827,32);
				when 3707 => sin_data_int <= to_signed(-562,32); cos_data_int <= to_signed(828,32);
				when 3708 => sin_data_int <= to_signed(-561,32); cos_data_int <= to_signed(829,32);
				when 3709 => sin_data_int <= to_signed(-559,32); cos_data_int <= to_signed(830,32);
				when 3710 => sin_data_int <= to_signed(-558,32); cos_data_int <= to_signed(831,32);
				when 3711 => sin_data_int <= to_signed(-557,32); cos_data_int <= to_signed(831,32);
				when 3712 => sin_data_int <= to_signed(-556,32); cos_data_int <= to_signed(832,32);
				when 3713 => sin_data_int <= to_signed(-554,32); cos_data_int <= to_signed(833,32);
				when 3714 => sin_data_int <= to_signed(-553,32); cos_data_int <= to_signed(834,32);
				when 3715 => sin_data_int <= to_signed(-552,32); cos_data_int <= to_signed(835,32);
				when 3716 => sin_data_int <= to_signed(-550,32); cos_data_int <= to_signed(836,32);
				when 3717 => sin_data_int <= to_signed(-549,32); cos_data_int <= to_signed(837,32);
				when 3718 => sin_data_int <= to_signed(-548,32); cos_data_int <= to_signed(837,32);
				when 3719 => sin_data_int <= to_signed(-547,32); cos_data_int <= to_signed(838,32);
				when 3720 => sin_data_int <= to_signed(-545,32); cos_data_int <= to_signed(839,32);
				when 3721 => sin_data_int <= to_signed(-544,32); cos_data_int <= to_signed(840,32);
				when 3722 => sin_data_int <= to_signed(-543,32); cos_data_int <= to_signed(841,32);
				when 3723 => sin_data_int <= to_signed(-541,32); cos_data_int <= to_signed(842,32);
				when 3724 => sin_data_int <= to_signed(-540,32); cos_data_int <= to_signed(842,32);
				when 3725 => sin_data_int <= to_signed(-539,32); cos_data_int <= to_signed(843,32);
				when 3726 => sin_data_int <= to_signed(-538,32); cos_data_int <= to_signed(844,32);
				when 3727 => sin_data_int <= to_signed(-536,32); cos_data_int <= to_signed(845,32);
				when 3728 => sin_data_int <= to_signed(-535,32); cos_data_int <= to_signed(846,32);
				when 3729 => sin_data_int <= to_signed(-534,32); cos_data_int <= to_signed(846,32);
				when 3730 => sin_data_int <= to_signed(-532,32); cos_data_int <= to_signed(847,32);
				when 3731 => sin_data_int <= to_signed(-531,32); cos_data_int <= to_signed(848,32);
				when 3732 => sin_data_int <= to_signed(-530,32); cos_data_int <= to_signed(849,32);
				when 3733 => sin_data_int <= to_signed(-529,32); cos_data_int <= to_signed(850,32);
				when 3734 => sin_data_int <= to_signed(-527,32); cos_data_int <= to_signed(851,32);
				when 3735 => sin_data_int <= to_signed(-526,32); cos_data_int <= to_signed(851,32);
				when 3736 => sin_data_int <= to_signed(-525,32); cos_data_int <= to_signed(852,32);
				when 3737 => sin_data_int <= to_signed(-523,32); cos_data_int <= to_signed(853,32);
				when 3738 => sin_data_int <= to_signed(-522,32); cos_data_int <= to_signed(854,32);
				when 3739 => sin_data_int <= to_signed(-521,32); cos_data_int <= to_signed(855,32);
				when 3740 => sin_data_int <= to_signed(-519,32); cos_data_int <= to_signed(855,32);
				when 3741 => sin_data_int <= to_signed(-518,32); cos_data_int <= to_signed(856,32);
				when 3742 => sin_data_int <= to_signed(-517,32); cos_data_int <= to_signed(857,32);
				when 3743 => sin_data_int <= to_signed(-515,32); cos_data_int <= to_signed(858,32);
				when 3744 => sin_data_int <= to_signed(-514,32); cos_data_int <= to_signed(859,32);
				when 3745 => sin_data_int <= to_signed(-513,32); cos_data_int <= to_signed(859,32);
				when 3746 => sin_data_int <= to_signed(-511,32); cos_data_int <= to_signed(860,32);
				when 3747 => sin_data_int <= to_signed(-510,32); cos_data_int <= to_signed(861,32);
				when 3748 => sin_data_int <= to_signed(-509,32); cos_data_int <= to_signed(862,32);
				when 3749 => sin_data_int <= to_signed(-508,32); cos_data_int <= to_signed(862,32);
				when 3750 => sin_data_int <= to_signed(-506,32); cos_data_int <= to_signed(863,32);
				when 3751 => sin_data_int <= to_signed(-505,32); cos_data_int <= to_signed(864,32);
				when 3752 => sin_data_int <= to_signed(-504,32); cos_data_int <= to_signed(865,32);
				when 3753 => sin_data_int <= to_signed(-502,32); cos_data_int <= to_signed(866,32);
				when 3754 => sin_data_int <= to_signed(-501,32); cos_data_int <= to_signed(866,32);
				when 3755 => sin_data_int <= to_signed(-500,32); cos_data_int <= to_signed(867,32);
				when 3756 => sin_data_int <= to_signed(-498,32); cos_data_int <= to_signed(868,32);
				when 3757 => sin_data_int <= to_signed(-497,32); cos_data_int <= to_signed(869,32);
				when 3758 => sin_data_int <= to_signed(-496,32); cos_data_int <= to_signed(869,32);
				when 3759 => sin_data_int <= to_signed(-494,32); cos_data_int <= to_signed(870,32);
				when 3760 => sin_data_int <= to_signed(-493,32); cos_data_int <= to_signed(871,32);
				when 3761 => sin_data_int <= to_signed(-492,32); cos_data_int <= to_signed(872,32);
				when 3762 => sin_data_int <= to_signed(-490,32); cos_data_int <= to_signed(872,32);
				when 3763 => sin_data_int <= to_signed(-489,32); cos_data_int <= to_signed(873,32);
				when 3764 => sin_data_int <= to_signed(-488,32); cos_data_int <= to_signed(874,32);
				when 3765 => sin_data_int <= to_signed(-486,32); cos_data_int <= to_signed(875,32);
				when 3766 => sin_data_int <= to_signed(-485,32); cos_data_int <= to_signed(875,32);
				when 3767 => sin_data_int <= to_signed(-484,32); cos_data_int <= to_signed(876,32);
				when 3768 => sin_data_int <= to_signed(-482,32); cos_data_int <= to_signed(877,32);
				when 3769 => sin_data_int <= to_signed(-481,32); cos_data_int <= to_signed(878,32);
				when 3770 => sin_data_int <= to_signed(-479,32); cos_data_int <= to_signed(878,32);
				when 3771 => sin_data_int <= to_signed(-478,32); cos_data_int <= to_signed(879,32);
				when 3772 => sin_data_int <= to_signed(-477,32); cos_data_int <= to_signed(880,32);
				when 3773 => sin_data_int <= to_signed(-475,32); cos_data_int <= to_signed(880,32);
				when 3774 => sin_data_int <= to_signed(-474,32); cos_data_int <= to_signed(881,32);
				when 3775 => sin_data_int <= to_signed(-473,32); cos_data_int <= to_signed(882,32);
				when 3776 => sin_data_int <= to_signed(-471,32); cos_data_int <= to_signed(883,32);
				when 3777 => sin_data_int <= to_signed(-470,32); cos_data_int <= to_signed(883,32);
				when 3778 => sin_data_int <= to_signed(-469,32); cos_data_int <= to_signed(884,32);
				when 3779 => sin_data_int <= to_signed(-467,32); cos_data_int <= to_signed(885,32);
				when 3780 => sin_data_int <= to_signed(-466,32); cos_data_int <= to_signed(886,32);
				when 3781 => sin_data_int <= to_signed(-465,32); cos_data_int <= to_signed(886,32);
				when 3782 => sin_data_int <= to_signed(-463,32); cos_data_int <= to_signed(887,32);
				when 3783 => sin_data_int <= to_signed(-462,32); cos_data_int <= to_signed(888,32);
				when 3784 => sin_data_int <= to_signed(-461,32); cos_data_int <= to_signed(888,32);
				when 3785 => sin_data_int <= to_signed(-459,32); cos_data_int <= to_signed(889,32);
				when 3786 => sin_data_int <= to_signed(-458,32); cos_data_int <= to_signed(890,32);
				when 3787 => sin_data_int <= to_signed(-456,32); cos_data_int <= to_signed(890,32);
				when 3788 => sin_data_int <= to_signed(-455,32); cos_data_int <= to_signed(891,32);
				when 3789 => sin_data_int <= to_signed(-454,32); cos_data_int <= to_signed(892,32);
				when 3790 => sin_data_int <= to_signed(-452,32); cos_data_int <= to_signed(893,32);
				when 3791 => sin_data_int <= to_signed(-451,32); cos_data_int <= to_signed(893,32);
				when 3792 => sin_data_int <= to_signed(-450,32); cos_data_int <= to_signed(894,32);
				when 3793 => sin_data_int <= to_signed(-448,32); cos_data_int <= to_signed(895,32);
				when 3794 => sin_data_int <= to_signed(-447,32); cos_data_int <= to_signed(895,32);
				when 3795 => sin_data_int <= to_signed(-445,32); cos_data_int <= to_signed(896,32);
				when 3796 => sin_data_int <= to_signed(-444,32); cos_data_int <= to_signed(897,32);
				when 3797 => sin_data_int <= to_signed(-443,32); cos_data_int <= to_signed(897,32);
				when 3798 => sin_data_int <= to_signed(-441,32); cos_data_int <= to_signed(898,32);
				when 3799 => sin_data_int <= to_signed(-440,32); cos_data_int <= to_signed(899,32);
				when 3800 => sin_data_int <= to_signed(-439,32); cos_data_int <= to_signed(899,32);
				when 3801 => sin_data_int <= to_signed(-437,32); cos_data_int <= to_signed(900,32);
				when 3802 => sin_data_int <= to_signed(-436,32); cos_data_int <= to_signed(901,32);
				when 3803 => sin_data_int <= to_signed(-434,32); cos_data_int <= to_signed(901,32);
				when 3804 => sin_data_int <= to_signed(-433,32); cos_data_int <= to_signed(902,32);
				when 3805 => sin_data_int <= to_signed(-432,32); cos_data_int <= to_signed(903,32);
				when 3806 => sin_data_int <= to_signed(-430,32); cos_data_int <= to_signed(903,32);
				when 3807 => sin_data_int <= to_signed(-429,32); cos_data_int <= to_signed(904,32);
				when 3808 => sin_data_int <= to_signed(-428,32); cos_data_int <= to_signed(905,32);
				when 3809 => sin_data_int <= to_signed(-426,32); cos_data_int <= to_signed(905,32);
				when 3810 => sin_data_int <= to_signed(-425,32); cos_data_int <= to_signed(906,32);
				when 3811 => sin_data_int <= to_signed(-423,32); cos_data_int <= to_signed(907,32);
				when 3812 => sin_data_int <= to_signed(-422,32); cos_data_int <= to_signed(907,32);
				when 3813 => sin_data_int <= to_signed(-421,32); cos_data_int <= to_signed(908,32);
				when 3814 => sin_data_int <= to_signed(-419,32); cos_data_int <= to_signed(909,32);
				when 3815 => sin_data_int <= to_signed(-418,32); cos_data_int <= to_signed(909,32);
				when 3816 => sin_data_int <= to_signed(-416,32); cos_data_int <= to_signed(910,32);
				when 3817 => sin_data_int <= to_signed(-415,32); cos_data_int <= to_signed(910,32);
				when 3818 => sin_data_int <= to_signed(-414,32); cos_data_int <= to_signed(911,32);
				when 3819 => sin_data_int <= to_signed(-412,32); cos_data_int <= to_signed(912,32);
				when 3820 => sin_data_int <= to_signed(-411,32); cos_data_int <= to_signed(912,32);
				when 3821 => sin_data_int <= to_signed(-409,32); cos_data_int <= to_signed(913,32);
				when 3822 => sin_data_int <= to_signed(-408,32); cos_data_int <= to_signed(914,32);
				when 3823 => sin_data_int <= to_signed(-407,32); cos_data_int <= to_signed(914,32);
				when 3824 => sin_data_int <= to_signed(-405,32); cos_data_int <= to_signed(915,32);
				when 3825 => sin_data_int <= to_signed(-404,32); cos_data_int <= to_signed(915,32);
				when 3826 => sin_data_int <= to_signed(-402,32); cos_data_int <= to_signed(916,32);
				when 3827 => sin_data_int <= to_signed(-401,32); cos_data_int <= to_signed(917,32);
				when 3828 => sin_data_int <= to_signed(-400,32); cos_data_int <= to_signed(917,32);
				when 3829 => sin_data_int <= to_signed(-398,32); cos_data_int <= to_signed(918,32);
				when 3830 => sin_data_int <= to_signed(-397,32); cos_data_int <= to_signed(919,32);
				when 3831 => sin_data_int <= to_signed(-395,32); cos_data_int <= to_signed(919,32);
				when 3832 => sin_data_int <= to_signed(-394,32); cos_data_int <= to_signed(920,32);
				when 3833 => sin_data_int <= to_signed(-393,32); cos_data_int <= to_signed(920,32);
				when 3834 => sin_data_int <= to_signed(-391,32); cos_data_int <= to_signed(921,32);
				when 3835 => sin_data_int <= to_signed(-390,32); cos_data_int <= to_signed(922,32);
				when 3836 => sin_data_int <= to_signed(-388,32); cos_data_int <= to_signed(922,32);
				when 3837 => sin_data_int <= to_signed(-387,32); cos_data_int <= to_signed(923,32);
				when 3838 => sin_data_int <= to_signed(-386,32); cos_data_int <= to_signed(923,32);
				when 3839 => sin_data_int <= to_signed(-384,32); cos_data_int <= to_signed(924,32);
				when 3840 => sin_data_int <= to_signed(-383,32); cos_data_int <= to_signed(924,32);
				when 3841 => sin_data_int <= to_signed(-381,32); cos_data_int <= to_signed(925,32);
				when 3842 => sin_data_int <= to_signed(-380,32); cos_data_int <= to_signed(926,32);
				when 3843 => sin_data_int <= to_signed(-378,32); cos_data_int <= to_signed(926,32);
				when 3844 => sin_data_int <= to_signed(-377,32); cos_data_int <= to_signed(927,32);
				when 3845 => sin_data_int <= to_signed(-376,32); cos_data_int <= to_signed(927,32);
				when 3846 => sin_data_int <= to_signed(-374,32); cos_data_int <= to_signed(928,32);
				when 3847 => sin_data_int <= to_signed(-373,32); cos_data_int <= to_signed(929,32);
				when 3848 => sin_data_int <= to_signed(-371,32); cos_data_int <= to_signed(929,32);
				when 3849 => sin_data_int <= to_signed(-370,32); cos_data_int <= to_signed(930,32);
				when 3850 => sin_data_int <= to_signed(-368,32); cos_data_int <= to_signed(930,32);
				when 3851 => sin_data_int <= to_signed(-367,32); cos_data_int <= to_signed(931,32);
				when 3852 => sin_data_int <= to_signed(-366,32); cos_data_int <= to_signed(931,32);
				when 3853 => sin_data_int <= to_signed(-364,32); cos_data_int <= to_signed(932,32);
				when 3854 => sin_data_int <= to_signed(-363,32); cos_data_int <= to_signed(932,32);
				when 3855 => sin_data_int <= to_signed(-361,32); cos_data_int <= to_signed(933,32);
				when 3856 => sin_data_int <= to_signed(-360,32); cos_data_int <= to_signed(934,32);
				when 3857 => sin_data_int <= to_signed(-358,32); cos_data_int <= to_signed(934,32);
				when 3858 => sin_data_int <= to_signed(-357,32); cos_data_int <= to_signed(935,32);
				when 3859 => sin_data_int <= to_signed(-356,32); cos_data_int <= to_signed(935,32);
				when 3860 => sin_data_int <= to_signed(-354,32); cos_data_int <= to_signed(936,32);
				when 3861 => sin_data_int <= to_signed(-353,32); cos_data_int <= to_signed(936,32);
				when 3862 => sin_data_int <= to_signed(-351,32); cos_data_int <= to_signed(937,32);
				when 3863 => sin_data_int <= to_signed(-350,32); cos_data_int <= to_signed(937,32);
				when 3864 => sin_data_int <= to_signed(-348,32); cos_data_int <= to_signed(938,32);
				when 3865 => sin_data_int <= to_signed(-347,32); cos_data_int <= to_signed(938,32);
				when 3866 => sin_data_int <= to_signed(-346,32); cos_data_int <= to_signed(939,32);
				when 3867 => sin_data_int <= to_signed(-344,32); cos_data_int <= to_signed(939,32);
				when 3868 => sin_data_int <= to_signed(-343,32); cos_data_int <= to_signed(940,32);
				when 3869 => sin_data_int <= to_signed(-341,32); cos_data_int <= to_signed(941,32);
				when 3870 => sin_data_int <= to_signed(-340,32); cos_data_int <= to_signed(941,32);
				when 3871 => sin_data_int <= to_signed(-338,32); cos_data_int <= to_signed(942,32);
				when 3872 => sin_data_int <= to_signed(-337,32); cos_data_int <= to_signed(942,32);
				when 3873 => sin_data_int <= to_signed(-335,32); cos_data_int <= to_signed(943,32);
				when 3874 => sin_data_int <= to_signed(-334,32); cos_data_int <= to_signed(943,32);
				when 3875 => sin_data_int <= to_signed(-333,32); cos_data_int <= to_signed(944,32);
				when 3876 => sin_data_int <= to_signed(-331,32); cos_data_int <= to_signed(944,32);
				when 3877 => sin_data_int <= to_signed(-330,32); cos_data_int <= to_signed(945,32);
				when 3878 => sin_data_int <= to_signed(-328,32); cos_data_int <= to_signed(945,32);
				when 3879 => sin_data_int <= to_signed(-327,32); cos_data_int <= to_signed(946,32);
				when 3880 => sin_data_int <= to_signed(-325,32); cos_data_int <= to_signed(946,32);
				when 3881 => sin_data_int <= to_signed(-324,32); cos_data_int <= to_signed(947,32);
				when 3882 => sin_data_int <= to_signed(-322,32); cos_data_int <= to_signed(947,32);
				when 3883 => sin_data_int <= to_signed(-321,32); cos_data_int <= to_signed(948,32);
				when 3884 => sin_data_int <= to_signed(-320,32); cos_data_int <= to_signed(948,32);
				when 3885 => sin_data_int <= to_signed(-318,32); cos_data_int <= to_signed(949,32);
				when 3886 => sin_data_int <= to_signed(-317,32); cos_data_int <= to_signed(949,32);
				when 3887 => sin_data_int <= to_signed(-315,32); cos_data_int <= to_signed(950,32);
				when 3888 => sin_data_int <= to_signed(-314,32); cos_data_int <= to_signed(950,32);
				when 3889 => sin_data_int <= to_signed(-312,32); cos_data_int <= to_signed(950,32);
				when 3890 => sin_data_int <= to_signed(-311,32); cos_data_int <= to_signed(951,32);
				when 3891 => sin_data_int <= to_signed(-309,32); cos_data_int <= to_signed(951,32);
				when 3892 => sin_data_int <= to_signed(-308,32); cos_data_int <= to_signed(952,32);
				when 3893 => sin_data_int <= to_signed(-306,32); cos_data_int <= to_signed(952,32);
				when 3894 => sin_data_int <= to_signed(-305,32); cos_data_int <= to_signed(953,32);
				when 3895 => sin_data_int <= to_signed(-303,32); cos_data_int <= to_signed(953,32);
				when 3896 => sin_data_int <= to_signed(-302,32); cos_data_int <= to_signed(954,32);
				when 3897 => sin_data_int <= to_signed(-301,32); cos_data_int <= to_signed(954,32);
				when 3898 => sin_data_int <= to_signed(-299,32); cos_data_int <= to_signed(955,32);
				when 3899 => sin_data_int <= to_signed(-298,32); cos_data_int <= to_signed(955,32);
				when 3900 => sin_data_int <= to_signed(-296,32); cos_data_int <= to_signed(956,32);
				when 3901 => sin_data_int <= to_signed(-295,32); cos_data_int <= to_signed(956,32);
				when 3902 => sin_data_int <= to_signed(-293,32); cos_data_int <= to_signed(956,32);
				when 3903 => sin_data_int <= to_signed(-292,32); cos_data_int <= to_signed(957,32);
				when 3904 => sin_data_int <= to_signed(-290,32); cos_data_int <= to_signed(957,32);
				when 3905 => sin_data_int <= to_signed(-289,32); cos_data_int <= to_signed(958,32);
				when 3906 => sin_data_int <= to_signed(-287,32); cos_data_int <= to_signed(958,32);
				when 3907 => sin_data_int <= to_signed(-286,32); cos_data_int <= to_signed(959,32);
				when 3908 => sin_data_int <= to_signed(-284,32); cos_data_int <= to_signed(959,32);
				when 3909 => sin_data_int <= to_signed(-283,32); cos_data_int <= to_signed(960,32);
				when 3910 => sin_data_int <= to_signed(-281,32); cos_data_int <= to_signed(960,32);
				when 3911 => sin_data_int <= to_signed(-280,32); cos_data_int <= to_signed(960,32);
				when 3912 => sin_data_int <= to_signed(-279,32); cos_data_int <= to_signed(961,32);
				when 3913 => sin_data_int <= to_signed(-277,32); cos_data_int <= to_signed(961,32);
				when 3914 => sin_data_int <= to_signed(-276,32); cos_data_int <= to_signed(962,32);
				when 3915 => sin_data_int <= to_signed(-274,32); cos_data_int <= to_signed(962,32);
				when 3916 => sin_data_int <= to_signed(-273,32); cos_data_int <= to_signed(963,32);
				when 3917 => sin_data_int <= to_signed(-271,32); cos_data_int <= to_signed(963,32);
				when 3918 => sin_data_int <= to_signed(-270,32); cos_data_int <= to_signed(963,32);
				when 3919 => sin_data_int <= to_signed(-268,32); cos_data_int <= to_signed(964,32);
				when 3920 => sin_data_int <= to_signed(-267,32); cos_data_int <= to_signed(964,32);
				when 3921 => sin_data_int <= to_signed(-265,32); cos_data_int <= to_signed(965,32);
				when 3922 => sin_data_int <= to_signed(-264,32); cos_data_int <= to_signed(965,32);
				when 3923 => sin_data_int <= to_signed(-262,32); cos_data_int <= to_signed(965,32);
				when 3924 => sin_data_int <= to_signed(-261,32); cos_data_int <= to_signed(966,32);
				when 3925 => sin_data_int <= to_signed(-259,32); cos_data_int <= to_signed(966,32);
				when 3926 => sin_data_int <= to_signed(-258,32); cos_data_int <= to_signed(967,32);
				when 3927 => sin_data_int <= to_signed(-256,32); cos_data_int <= to_signed(967,32);
				when 3928 => sin_data_int <= to_signed(-255,32); cos_data_int <= to_signed(967,32);
				when 3929 => sin_data_int <= to_signed(-253,32); cos_data_int <= to_signed(968,32);
				when 3930 => sin_data_int <= to_signed(-252,32); cos_data_int <= to_signed(968,32);
				when 3931 => sin_data_int <= to_signed(-250,32); cos_data_int <= to_signed(969,32);
				when 3932 => sin_data_int <= to_signed(-249,32); cos_data_int <= to_signed(969,32);
				when 3933 => sin_data_int <= to_signed(-247,32); cos_data_int <= to_signed(969,32);
				when 3934 => sin_data_int <= to_signed(-246,32); cos_data_int <= to_signed(970,32);
				when 3935 => sin_data_int <= to_signed(-244,32); cos_data_int <= to_signed(970,32);
				when 3936 => sin_data_int <= to_signed(-243,32); cos_data_int <= to_signed(970,32);
				when 3937 => sin_data_int <= to_signed(-241,32); cos_data_int <= to_signed(971,32);
				when 3938 => sin_data_int <= to_signed(-240,32); cos_data_int <= to_signed(971,32);
				when 3939 => sin_data_int <= to_signed(-239,32); cos_data_int <= to_signed(972,32);
				when 3940 => sin_data_int <= to_signed(-237,32); cos_data_int <= to_signed(972,32);
				when 3941 => sin_data_int <= to_signed(-236,32); cos_data_int <= to_signed(972,32);
				when 3942 => sin_data_int <= to_signed(-234,32); cos_data_int <= to_signed(973,32);
				when 3943 => sin_data_int <= to_signed(-233,32); cos_data_int <= to_signed(973,32);
				when 3944 => sin_data_int <= to_signed(-231,32); cos_data_int <= to_signed(973,32);
				when 3945 => sin_data_int <= to_signed(-230,32); cos_data_int <= to_signed(974,32);
				when 3946 => sin_data_int <= to_signed(-228,32); cos_data_int <= to_signed(974,32);
				when 3947 => sin_data_int <= to_signed(-227,32); cos_data_int <= to_signed(974,32);
				when 3948 => sin_data_int <= to_signed(-225,32); cos_data_int <= to_signed(975,32);
				when 3949 => sin_data_int <= to_signed(-224,32); cos_data_int <= to_signed(975,32);
				when 3950 => sin_data_int <= to_signed(-222,32); cos_data_int <= to_signed(975,32);
				when 3951 => sin_data_int <= to_signed(-221,32); cos_data_int <= to_signed(976,32);
				when 3952 => sin_data_int <= to_signed(-219,32); cos_data_int <= to_signed(976,32);
				when 3953 => sin_data_int <= to_signed(-218,32); cos_data_int <= to_signed(976,32);
				when 3954 => sin_data_int <= to_signed(-216,32); cos_data_int <= to_signed(977,32);
				when 3955 => sin_data_int <= to_signed(-215,32); cos_data_int <= to_signed(977,32);
				when 3956 => sin_data_int <= to_signed(-213,32); cos_data_int <= to_signed(977,32);
				when 3957 => sin_data_int <= to_signed(-212,32); cos_data_int <= to_signed(978,32);
				when 3958 => sin_data_int <= to_signed(-210,32); cos_data_int <= to_signed(978,32);
				when 3959 => sin_data_int <= to_signed(-209,32); cos_data_int <= to_signed(978,32);
				when 3960 => sin_data_int <= to_signed(-207,32); cos_data_int <= to_signed(979,32);
				when 3961 => sin_data_int <= to_signed(-206,32); cos_data_int <= to_signed(979,32);
				when 3962 => sin_data_int <= to_signed(-204,32); cos_data_int <= to_signed(979,32);
				when 3963 => sin_data_int <= to_signed(-203,32); cos_data_int <= to_signed(980,32);
				when 3964 => sin_data_int <= to_signed(-201,32); cos_data_int <= to_signed(980,32);
				when 3965 => sin_data_int <= to_signed(-200,32); cos_data_int <= to_signed(980,32);
				when 3966 => sin_data_int <= to_signed(-198,32); cos_data_int <= to_signed(980,32);
				when 3967 => sin_data_int <= to_signed(-197,32); cos_data_int <= to_signed(981,32);
				when 3968 => sin_data_int <= to_signed(-195,32); cos_data_int <= to_signed(981,32);
				when 3969 => sin_data_int <= to_signed(-194,32); cos_data_int <= to_signed(981,32);
				when 3970 => sin_data_int <= to_signed(-192,32); cos_data_int <= to_signed(982,32);
				when 3971 => sin_data_int <= to_signed(-191,32); cos_data_int <= to_signed(982,32);
				when 3972 => sin_data_int <= to_signed(-189,32); cos_data_int <= to_signed(982,32);
				when 3973 => sin_data_int <= to_signed(-188,32); cos_data_int <= to_signed(983,32);
				when 3974 => sin_data_int <= to_signed(-186,32); cos_data_int <= to_signed(983,32);
				when 3975 => sin_data_int <= to_signed(-185,32); cos_data_int <= to_signed(983,32);
				when 3976 => sin_data_int <= to_signed(-183,32); cos_data_int <= to_signed(983,32);
				when 3977 => sin_data_int <= to_signed(-182,32); cos_data_int <= to_signed(984,32);
				when 3978 => sin_data_int <= to_signed(-180,32); cos_data_int <= to_signed(984,32);
				when 3979 => sin_data_int <= to_signed(-179,32); cos_data_int <= to_signed(984,32);
				when 3980 => sin_data_int <= to_signed(-177,32); cos_data_int <= to_signed(984,32);
				when 3981 => sin_data_int <= to_signed(-175,32); cos_data_int <= to_signed(985,32);
				when 3982 => sin_data_int <= to_signed(-174,32); cos_data_int <= to_signed(985,32);
				when 3983 => sin_data_int <= to_signed(-172,32); cos_data_int <= to_signed(985,32);
				when 3984 => sin_data_int <= to_signed(-171,32); cos_data_int <= to_signed(986,32);
				when 3985 => sin_data_int <= to_signed(-169,32); cos_data_int <= to_signed(986,32);
				when 3986 => sin_data_int <= to_signed(-168,32); cos_data_int <= to_signed(986,32);
				when 3987 => sin_data_int <= to_signed(-166,32); cos_data_int <= to_signed(986,32);
				when 3988 => sin_data_int <= to_signed(-165,32); cos_data_int <= to_signed(987,32);
				when 3989 => sin_data_int <= to_signed(-163,32); cos_data_int <= to_signed(987,32);
				when 3990 => sin_data_int <= to_signed(-162,32); cos_data_int <= to_signed(987,32);
				when 3991 => sin_data_int <= to_signed(-160,32); cos_data_int <= to_signed(987,32);
				when 3992 => sin_data_int <= to_signed(-159,32); cos_data_int <= to_signed(988,32);
				when 3993 => sin_data_int <= to_signed(-157,32); cos_data_int <= to_signed(988,32);
				when 3994 => sin_data_int <= to_signed(-156,32); cos_data_int <= to_signed(988,32);
				when 3995 => sin_data_int <= to_signed(-154,32); cos_data_int <= to_signed(988,32);
				when 3996 => sin_data_int <= to_signed(-153,32); cos_data_int <= to_signed(988,32);
				when 3997 => sin_data_int <= to_signed(-151,32); cos_data_int <= to_signed(989,32);
				when 3998 => sin_data_int <= to_signed(-150,32); cos_data_int <= to_signed(989,32);
				when 3999 => sin_data_int <= to_signed(-148,32); cos_data_int <= to_signed(989,32);
				when 4000 => sin_data_int <= to_signed(-147,32); cos_data_int <= to_signed(989,32);
				when 4001 => sin_data_int <= to_signed(-145,32); cos_data_int <= to_signed(990,32);
				when 4002 => sin_data_int <= to_signed(-144,32); cos_data_int <= to_signed(990,32);
				when 4003 => sin_data_int <= to_signed(-142,32); cos_data_int <= to_signed(990,32);
				when 4004 => sin_data_int <= to_signed(-141,32); cos_data_int <= to_signed(990,32);
				when 4005 => sin_data_int <= to_signed(-139,32); cos_data_int <= to_signed(990,32);
				when 4006 => sin_data_int <= to_signed(-138,32); cos_data_int <= to_signed(991,32);
				when 4007 => sin_data_int <= to_signed(-136,32); cos_data_int <= to_signed(991,32);
				when 4008 => sin_data_int <= to_signed(-135,32); cos_data_int <= to_signed(991,32);
				when 4009 => sin_data_int <= to_signed(-133,32); cos_data_int <= to_signed(991,32);
				when 4010 => sin_data_int <= to_signed(-132,32); cos_data_int <= to_signed(992,32);
				when 4011 => sin_data_int <= to_signed(-130,32); cos_data_int <= to_signed(992,32);
				when 4012 => sin_data_int <= to_signed(-128,32); cos_data_int <= to_signed(992,32);
				when 4013 => sin_data_int <= to_signed(-127,32); cos_data_int <= to_signed(992,32);
				when 4014 => sin_data_int <= to_signed(-125,32); cos_data_int <= to_signed(992,32);
				when 4015 => sin_data_int <= to_signed(-124,32); cos_data_int <= to_signed(992,32);
				when 4016 => sin_data_int <= to_signed(-122,32); cos_data_int <= to_signed(993,32);
				when 4017 => sin_data_int <= to_signed(-121,32); cos_data_int <= to_signed(993,32);
				when 4018 => sin_data_int <= to_signed(-119,32); cos_data_int <= to_signed(993,32);
				when 4019 => sin_data_int <= to_signed(-118,32); cos_data_int <= to_signed(993,32);
				when 4020 => sin_data_int <= to_signed(-116,32); cos_data_int <= to_signed(993,32);
				when 4021 => sin_data_int <= to_signed(-115,32); cos_data_int <= to_signed(994,32);
				when 4022 => sin_data_int <= to_signed(-113,32); cos_data_int <= to_signed(994,32);
				when 4023 => sin_data_int <= to_signed(-112,32); cos_data_int <= to_signed(994,32);
				when 4024 => sin_data_int <= to_signed(-110,32); cos_data_int <= to_signed(994,32);
				when 4025 => sin_data_int <= to_signed(-109,32); cos_data_int <= to_signed(994,32);
				when 4026 => sin_data_int <= to_signed(-107,32); cos_data_int <= to_signed(994,32);
				when 4027 => sin_data_int <= to_signed(-106,32); cos_data_int <= to_signed(995,32);
				when 4028 => sin_data_int <= to_signed(-104,32); cos_data_int <= to_signed(995,32);
				when 4029 => sin_data_int <= to_signed(-103,32); cos_data_int <= to_signed(995,32);
				when 4030 => sin_data_int <= to_signed(-101,32); cos_data_int <= to_signed(995,32);
				when 4031 => sin_data_int <= to_signed(-100,32); cos_data_int <= to_signed(995,32);
				when 4032 => sin_data_int <= to_signed(-98,32); cos_data_int <= to_signed(995,32);
				when 4033 => sin_data_int <= to_signed(-96,32); cos_data_int <= to_signed(995,32);
				when 4034 => sin_data_int <= to_signed(-95,32); cos_data_int <= to_signed(996,32);
				when 4035 => sin_data_int <= to_signed(-93,32); cos_data_int <= to_signed(996,32);
				when 4036 => sin_data_int <= to_signed(-92,32); cos_data_int <= to_signed(996,32);
				when 4037 => sin_data_int <= to_signed(-90,32); cos_data_int <= to_signed(996,32);
				when 4038 => sin_data_int <= to_signed(-89,32); cos_data_int <= to_signed(996,32);
				when 4039 => sin_data_int <= to_signed(-87,32); cos_data_int <= to_signed(996,32);
				when 4040 => sin_data_int <= to_signed(-86,32); cos_data_int <= to_signed(996,32);
				when 4041 => sin_data_int <= to_signed(-84,32); cos_data_int <= to_signed(997,32);
				when 4042 => sin_data_int <= to_signed(-83,32); cos_data_int <= to_signed(997,32);
				when 4043 => sin_data_int <= to_signed(-81,32); cos_data_int <= to_signed(997,32);
				when 4044 => sin_data_int <= to_signed(-80,32); cos_data_int <= to_signed(997,32);
				when 4045 => sin_data_int <= to_signed(-78,32); cos_data_int <= to_signed(997,32);
				when 4046 => sin_data_int <= to_signed(-77,32); cos_data_int <= to_signed(997,32);
				when 4047 => sin_data_int <= to_signed(-75,32); cos_data_int <= to_signed(997,32);
				when 4048 => sin_data_int <= to_signed(-74,32); cos_data_int <= to_signed(997,32);
				when 4049 => sin_data_int <= to_signed(-72,32); cos_data_int <= to_signed(998,32);
				when 4050 => sin_data_int <= to_signed(-71,32); cos_data_int <= to_signed(998,32);
				when 4051 => sin_data_int <= to_signed(-69,32); cos_data_int <= to_signed(998,32);
				when 4052 => sin_data_int <= to_signed(-67,32); cos_data_int <= to_signed(998,32);
				when 4053 => sin_data_int <= to_signed(-66,32); cos_data_int <= to_signed(998,32);
				when 4054 => sin_data_int <= to_signed(-64,32); cos_data_int <= to_signed(998,32);
				when 4055 => sin_data_int <= to_signed(-63,32); cos_data_int <= to_signed(998,32);
				when 4056 => sin_data_int <= to_signed(-61,32); cos_data_int <= to_signed(998,32);
				when 4057 => sin_data_int <= to_signed(-60,32); cos_data_int <= to_signed(998,32);
				when 4058 => sin_data_int <= to_signed(-58,32); cos_data_int <= to_signed(998,32);
				when 4059 => sin_data_int <= to_signed(-57,32); cos_data_int <= to_signed(998,32);
				when 4060 => sin_data_int <= to_signed(-55,32); cos_data_int <= to_signed(999,32);
				when 4061 => sin_data_int <= to_signed(-54,32); cos_data_int <= to_signed(999,32);
				when 4062 => sin_data_int <= to_signed(-52,32); cos_data_int <= to_signed(999,32);
				when 4063 => sin_data_int <= to_signed(-51,32); cos_data_int <= to_signed(999,32);
				when 4064 => sin_data_int <= to_signed(-49,32); cos_data_int <= to_signed(999,32);
				when 4065 => sin_data_int <= to_signed(-48,32); cos_data_int <= to_signed(999,32);
				when 4066 => sin_data_int <= to_signed(-46,32); cos_data_int <= to_signed(999,32);
				when 4067 => sin_data_int <= to_signed(-44,32); cos_data_int <= to_signed(999,32);
				when 4068 => sin_data_int <= to_signed(-43,32); cos_data_int <= to_signed(999,32);
				when 4069 => sin_data_int <= to_signed(-41,32); cos_data_int <= to_signed(999,32);
				when 4070 => sin_data_int <= to_signed(-40,32); cos_data_int <= to_signed(999,32);
				when 4071 => sin_data_int <= to_signed(-38,32); cos_data_int <= to_signed(999,32);
				when 4072 => sin_data_int <= to_signed(-37,32); cos_data_int <= to_signed(999,32);
				when 4073 => sin_data_int <= to_signed(-35,32); cos_data_int <= to_signed(999,32);
				when 4074 => sin_data_int <= to_signed(-34,32); cos_data_int <= to_signed(999,32);
				when 4075 => sin_data_int <= to_signed(-32,32); cos_data_int <= to_signed(1000,32);
				when 4076 => sin_data_int <= to_signed(-31,32); cos_data_int <= to_signed(1000,32);
				when 4077 => sin_data_int <= to_signed(-29,32); cos_data_int <= to_signed(1000,32);
				when 4078 => sin_data_int <= to_signed(-28,32); cos_data_int <= to_signed(1000,32);
				when 4079 => sin_data_int <= to_signed(-26,32); cos_data_int <= to_signed(1000,32);
				when 4080 => sin_data_int <= to_signed(-25,32); cos_data_int <= to_signed(1000,32);
				when 4081 => sin_data_int <= to_signed(-23,32); cos_data_int <= to_signed(1000,32);
				when 4082 => sin_data_int <= to_signed(-21,32); cos_data_int <= to_signed(1000,32);
				when 4083 => sin_data_int <= to_signed(-20,32); cos_data_int <= to_signed(1000,32);
				when 4084 => sin_data_int <= to_signed(-18,32); cos_data_int <= to_signed(1000,32);
				when 4085 => sin_data_int <= to_signed(-17,32); cos_data_int <= to_signed(1000,32);
				when 4086 => sin_data_int <= to_signed(-15,32); cos_data_int <= to_signed(1000,32);
				when 4087 => sin_data_int <= to_signed(-14,32); cos_data_int <= to_signed(1000,32);
				when 4088 => sin_data_int <= to_signed(-12,32); cos_data_int <= to_signed(1000,32);
				when 4089 => sin_data_int <= to_signed(-11,32); cos_data_int <= to_signed(1000,32);
				when 4090 => sin_data_int <= to_signed(-9,32); cos_data_int <= to_signed(1000,32);
				when 4091 => sin_data_int <= to_signed(-8,32); cos_data_int <= to_signed(1000,32);
				when 4092 => sin_data_int <= to_signed(-6,32); cos_data_int <= to_signed(1000,32);
				when 4093 => sin_data_int <= to_signed(-5,32); cos_data_int <= to_signed(1000,32);
				when 4094 => sin_data_int <= to_signed(-3,32); cos_data_int <= to_signed(1000,32);
				when 4095 => sin_data_int <= to_signed(-2,32); cos_data_int <= to_signed(1000,32);
				--when 4096 => sin_data_int <= to_signed(0,32); cos_data_int <= to_signed(1000,32);
            when others       => null;

         end case;

      end if;
   end if;
end process;


end rtl;
